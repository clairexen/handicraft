module testbox_0(input A, B, output Y);
assign Y = 0;
endmodule
