// generated from the data at http://visual6502.org/JSSim/

module MOS6502(vss, rdy, clk1out, irq, nmi, sync, vcc, ab0, ab1, ab2, ab3, ab4, ab5, ab6, ab7, ab8, ab9, ab10, ab11,
		ab12, ab13, ab14, ab15, db7, db6, db5, db4, db3, db2, db1, db0, rw, clk0, so, clk2out, res);

input vss, vcc, irq, nmi, clk0, res, rdy, so;
inout db7, db6, db5, db4, db3, db2, db1, db0;

output clk1out, clk2out, sync, rw;
output ab0, ab1, ab2, ab3, ab4, ab5, ab6, ab7, ab8, ab9, ab10, ab11, ab12, ab13, ab14, ab15;

wire \op-T5-rts , x2, net2, net3, \op-T0-tay , net5, net6, net7, net8, net9;
wire net10, net11, net12, adh6, net14, net15, net16, net17, net18, net19;
wire net20, net21, \~(AxBxC)2 , net23, net24, net25, notir4, pchp4, \~ABL7 , net29;
wire net31, p0, \~pchp5 , net34, net35, net36, net37, net38, \~pclp4 , pipeT2out;
wire \dpc42_DL/ADH , net42, net43, pipeUNK05, pipeVectorA2, net46, net47, dpc30_ADHPCH, pch5, net50;
wire net51, adh1, \op-lsr/ror/dec/inc , dasb0, net55, pipeUNK34, net57, \op-T3-abs-idx , dpc13_ORS, \op-T3-ind-y ;
wire net61, net62, dor7, y0, \(AxB)4.~C34 , net66, RESP, notalu6, net69, net70;
wire net71, pclp5, pipeUNK27, net74, net75, \op-T0-dex , Pout6, C34, net79, net80;
wire s2, db1, net83, \op-T2-ind-x , x4, net86, net87, net88, rdy, net90;
wire net91, \~ABH3 , net93, net94, net95, alub3, dor0, x1, pipeUNK04, net100;
wire net101, net102, irq, net104, net105, net106, \~ABL1 , net108, net109, \A+B2 ;
wire net111, net112, \~pchp1 , \~pchp2 , y6, notidl0, \A+B7 , net118, net119, \op-T3 ;
wire adl6, net122, net123, \~pchp3 , \PD-n-0xx0xx0x , net126, net127, net128, dpc20_ADDSB06, net130;
wire \op-T0-pla , net132, net133, net134, net135, net136, net137, net138, net139, dpc27_SBADH;
wire pchp3, C45, \~(A+B)0 , \op-sta/cmp , net146, net147, ab9, net149, net150, pipeUNK39;
wire net152, \~ABL0 , net154, \~(A+B)1 , clock2, \op-T2-stack-access , notdor7, res, net160, net161;
wire a3, net163, \DC78.phi2 , net165, sb5, \op-T0-tax , net168, net169, pipeVectorA1, net171;
wire net172, \(AxB)6.~C56 , db5, net176, \~(AxB)7 , abl6, \op-T0-txa , net180, nots7, net182;
wire s1, noty3, net185, net186, notRnWprepad, net188, net189, net190, net191, net192;
wire \(AxB)2.~C12 , notir0, ab15, net196, pipeUNK37, net198, pipeUNK09, net200, net201, net202;
wire dpc29_0ADH17, \op-T2-ADL/ADD , pch7, \~alucout , net207, pclp4, pchp1, net210, ab3, net212;
wire net213, dpc19_ADDSB7, pipeUNK10, \DA-AB2 , \0/ADL0 , net218, \op-T2-mem-zp , net220, net221, notdor0;
wire net223, net224, net225, net226, net227, net228, dpc28_0ADH0, ab8, net231, net232;
wire net233, abl5, alub6, net236, net237, net238, net239, idl5, net241, net242;
wire net243, \op-ror , \op-T0-txs , net246, dpc33_PCHDB, notRdy0, net249, \~aluresult1 , net251, \~op-set-C ;
wire net253, net254, net255, net256, \op-T0-tya , \op-T2-idx-x-xy , \op-jsr , net260, net261, net262;
wire dasb5, \~NMIG , net265, net266, net267, ab0, net269, net270, \op-T0-jsr , net272;
wire \op-T2-abs-access , \~(AxBxC)3 , net275, notalu2, \~aluresult5 , net278, net279, net280, \op-T4-mem-abs-idx , net282;
wire dpc37_PCLDB, net284, \op-T2-zp/zp-idx , \op-T0-tay/ldy-not-idx , abh2, net288, \~ABH6 , net291, pch1, net293;
wire pipeUNK20, \~(AxB1).C01 , \~aluresult4 , \~NMIP , net298, net299, net300, \op-T+-cmp , \PD-xxx010x1 , \op-T0-bit ;
wire \~aluresult7 , y3, net306, net307, \~(AxB)4 , \op-T2-jmp-abs , net310, net311, net312, net313;
wire alu5, adh3, net316, net317, net318, net319, net320, net321, net322, net323;
wire \op-inc/nop , dpc1_SBY, net326, net327, ir0, net329, net330, alu6, net332, DC78;
wire net334, net335, \~A.B6 , ir6, pipeUNK08, net339, net340, \op-T4 , \x-op-T3-ind-y , net343;
wire net344, net345, net346, net347, p3, ab13, \~A.B3 , net351, \op-T4-brk , RnWstretched;
wire \op-T4-abs-idx , net355, net356, pipeVectorA0, net358, net359, net360, pd1, dpc14_SRS, net363;
wire \~ABL4 , \PD-0xx0xx0x , net366, net367, net368, pd4, \op-T5-brk , \~(AxBxC)0 , net372, net373;
wire net374, net375, abl1, pcl6, net378, \dpc36_~IPC , net380, net381, \op-T0-iny/dey , net383;
wire net384, net385, net386, net387, net388, net389, net390, idl7, net392, net393;
wire notalu0, net395, net396, net397, net398, ab11, net400, alu0, net402, \op-T0-ora ;
wire \~(A+B)4 , net405, net406, adh0, net408, net409, net410, notalucout, adl0, dpc40_ADLPCL;
wire net415, net416, net417, nots0, net419, net420, clk2out, abh3, net423, net424;
wire AxB1, net426, \~C56 , net428, \~ABH7 , \short-circuit-branch-add , net431, net432, net433, \op-rmw ;
wire ab4, net436, dpc10_ADLADD, dpc38_PCLADL, Pout3, net440, net441, net442, pipeUNK06, dor3;
wire net445, \op-T5-rti/rts , \x-op-T3-abs-idx , x6, pipephi2Reset0, dasb2, ab1, net452, net453, net454;
wire net455, pipeUNK40, net457, net458, net459, net460, \x-op-T4-ind-y , net462, net463, idl3;
wire \~~alucout , net466, net467, net468, net469, net470, net471, net472, net473, net474;
wire net475, net476, \~A.B5 , net478, net479, net480, pclp2, net482, adh5, net484;
wire notx4, \~(AxBxC)5 , \op-T2-brk , pclp0, abh7, net490, net491, \op-T4-ind-y , idb7, net494;
wire notalu3, net496, notidl5, net499, C56, net501, pch2, net503, net504, C12;
wire net506, net507, net508, net509, net510, net511, net512, net513, net514, net515;
wire \DA-AxB2 , \op-store , net518, net519, net520, net521, \op-ORS , net523, net524, net525;
wire net526, notdor1, \xx-op-T5-jsr , notidl7, alua5, net531, \~(AxBxC)7 , net533, dpc23_SBAC, \~pchp7 ;
wire \~pclp7 , \pipeT-SYNC , net538, sync, \pd4.clearIR , net541, net543, net544, net545, \op-shift ;
wire net547, net548, dpc11_SBADD, net550, net551, \op-T0-php/pha , net553, \pipe~T0 , \(AxB)0.~C0in , net556;
wire net557, vss, \~notRdy0.delay , \C78.phi2 , pipeUNK22, net562, net564, noty4, net566, abl7;
wire net568, net569, net570, net571, net572, y2, dpc15_ANDS, \op-T0-adc/sbc , notidl1, net577;
wire net578, \op-T3-jsr , net580, net581, net582, net583, pch3, net585, net586, net587;
wire net588, x5, net590, net591, \~C67 , net593, \op-T0-jmp , net595, pipeUNK23, net597;
wire net598, net599, net600, nots5, net602, net603, net604, net605, alu4, \op-T3-mem-abs ;
wire net608, net609, net610, net611, net612, net613, pipeUNK31, y5, net616, net617;
wire net618, net619, net620, net621, pcl5, \DA-C01 , net624, net625, \branch-back , p1;
wire net628, net629, net630, net631, net632, net633, net634, net635, net636, net637;
wire net638, \ADL/ABL , AxB3, net641, net642, net643, net644, net645, net646, net647;
wire net648, \~(A+B)3 , db3, \~(AxBxC)4 , pchp6, net653, dpc7_SS, pcl2, net656, vcc;
wire net658, net659, \op-T3-branch , net661, net662, net663, net664, \op-T0-ldy-mem , net666, \pd5.clearIR ;
wire \~ABH4 , net669, net670, net671, ab14, net673, net674, IRQP, net676, \op-T3-abs/idx/ind ;
wire net678, dasb6, net680, \~A.B2 , \op-T0-tsx , pipedpc28, adl3, pipeUNK28, \0/ADL1 , Pout0;
wire net688, net689, t4, \op-asl/rol , net692, \A+B0 , net694, net695, net696, notalu1;
wire net698, \~DA-ADD2 , net700, \~(AxB)2 , notir1, net703, alub2, net705, pipeT3out, \~ABL2 ;
wire net708, net709, cp1, net711, \op-T2-jsr , abh1, net714, net715, net716, net717;
wire net718, net719, net720, net721, \~aluresult6 , pclp3, net724, \dpc22_~DSA , net726, a4;
wire net728, pipeUNK36, notx6, \~pclp6 , net732, net733, net734, net735, ab5, a0;
wire net738, net739, \~aluresult2 , dpc31_PCHPCH, net742, net743, DBZ, net745, dor1, net747;
wire net748, \op-T2-php , \~pchp6 , nots2, net753, net754, net755, net756, net757, pd0;
wire net759, net760, net761, net762, net763, \op-jmp , alu7, net766, net767, \~ABH2 ;
wire net769, \notRdy0.delay , \branch-back.phi1 , net772, net773, net774, abh5, \op-T5-jsr , x7, ONEBYTE;
wire net779, \~pchp0 , net781, net782, net783, \op-T5-rti , net785, \op-T+-dex , \op-T0-sbc , \op-T2 ;
wire net789, net790, \op-push/pull , \~TWOCYCLE.phi1 , net793, net794, net795, net796, net797, net798;
wire net799, net800, dpc0_YSB, net802, \A+B6 , \op-T4-brk/jsr , net805, net806, net807, alurawcout;
wire \pd1.clearIR , net810, net811, net812, net813, net814, net815, net816, \~(AxB5).C45 , net818;
wire net819, \~pchp4 , \ADH/ABH , \op-T+-adc/sbc , notdor3, net824, \~ABL3 , net826, D1x1, nots3;
wire pd5, net830, net831, pipeUNK19, idb6, net834, net835, net836, net837, net838;
wire net839, \~op-branch-bit6 , \~A.B1 , net842, y7, net844, net845, net846, net847, pipeUNK33;
wire net849, net850, \~TWOCYCLE , net852, net853, net854, net855, net856, \op-rti/rts , a5;
wire dpc9_DBADD, \~(AxB3).C23 , net861, net862, \dpc43_DL/DB , net864, net865, net866, net867, \~pclp3 ;
wire net869, idl1, net871, alu1, notdor4, dpc6_SBS, net875, net876, net877, net878;
wire fetch, net880, net881, net882, net883, \~(AxB)3 , net885, net886, ab6, \~IRQP ;
wire net889, notx2, net891, idb4, notalu5, pd3, notir6, net896, net897, dpc39_PCLPCL;
wire pipeUNK18, pcl4, \~DA-ADD1 , net902, net903, \op-T3-mem-zp-idx , net905, net906, \~ABH1 , t5;
wire alucin, net911, net912, net913, net914, net916, net917, \A+B4 , net919, net920;
wire dpc17_SUMS, net922, net923, net924, \~op-store , RESG, net927, net928, net929, net930;
wire net931, \op-T2-php/pha , net933, \op-SRS , net935, net936, net937, aluvout, net939, pipeT5out;
wire net941, net942, cclk, net944, db2, net946, net947, pch4, net949, \op-T+-cpx/cpy-abs ;
wire net951, net952, \~(AxB)1 , net954, pd2, net956, \~aluresult0 , net958, net959, pipeUNK32;
wire net961, net962, net963, net964, \~(AxBxC)1 , net966, nnT2BR, net968, net969, net970;
wire t2, net972, net973, pipeUNK02, net975, pclp1, alub0, a2, net979, net980;
wire noty5, net982, net983, dpc12_0ADD, \op-T0-ldx/tax/tsx , net986, notx0, net988, y4, net990;
wire idb1, net992, net993, net994, net995, irline3, abh6, net998, net999, net1000;
wire sb7, net1002, \~C23 , net1004, db0, \op-implied , net1007, pipeUNK29, dasb1, net1010;
wire pipeUNK11, net1012, net1013, net1014, dpc21_ADDADL, net1016, notx5, net1018, \PD-xxxx10x0 , net1020;
wire \A+B1 , pcl1, C23, net1024, noty0, net1026, net1027, net1028, nots6, net1030;
wire \op-T3-stack/bit/jmp , NMIP, net1033, net1034, \~DBE , pipephi2Reset0x, net1037, net1038, net1039, net1040;
wire net1041, H1x1, net1043, net1044, net1045, net1046, net1047, \~op-branch-done , net1049, \x-op-push/pull ;
wire pipeUNK16, \x-op-jmp , net1053, net1054, net1055, net1056, \op-T2-abs , net1058, net1059, dpc25_SBDB;
wire net1061, \~ABH0 , \~A.B4 , nots1, net1065, idl2, net1067, dpc8_nDBADD, net1069, net1070;
wire \~aluresult3 , net1072, net1073, \op-T0-shift-right-a , net1075, net1076, clearIR, pipeUNK17, \~pclp2 , net1080;
wire net1081, net1082, net1083, \~(A+B)6 , net1085, \op-T2-pha , net1087, dor4, net1089, net1090;
wire net1091, net1092, net1093, net1094, net1095, abl0, net1097, s5, net1099, net1100;
wire net1101, \~pclp1 , net1103, pipeUNK42, net1105, net1106, net1107, idb0, net1109, \branch-forward.phi1 ;
wire net1111, ir4, net1113, \op-T0-clc/sec , net1115, idl6, net1117, net1118, Pout4, net1120;
wire net1121, \~C12 , notalu7, net1124, notir3, net1126, \~ABH5 , net1129, net1130, \pipe~WR.phi2 ;
wire net1132, net1133, \~VEC , net1135, a6, net1137, noty1, pcl0, net1140, net1141;
wire alua4, abh4, \DA-C45 , net1145, alucout, net1147, y1, net1149, sb1, net1151;
wire net1152, net1153, net1154, \x-op-T+-adc/sbc , rw, net1157, net1158, net1159, adh4, net1161;
wire net1162, clk1out, \op-clv , notalucin, net1166, alua0, \op-T5-ind-y , net1169, net1170, clk0;
wire net1172, \x-op-T0-tya , \~op-branch-bit7 , net1175, pipeUNK21, net1177, net1178, net1179, net1180, net1181;
wire notir2, net1183, net1184, \short-circuit-idx-add , dpc3_SBX, net1187, sb3, net1189, net1190, net1191;
wire net1192, \0/ADL2 , net1194, net1195, \op-SUMS , \~(AxBxC)6 , net1198, net1199, DBNeg, \dpc18_~DAA ;
wire net1202, net1203, \op-T2-ind-y , net1205, pchp7, net1209, \op-T5-ind-x , net1211, s6, net1213;
wire net1214, net1215, x0, \~(AxB7).C67 , net1218, net1219, AxB5, net1221, net1222, net1223;
wire net1224, net1225, \op-T0-plp , \~pclp0 , \op-ANDS , net1229, net1230, net1231, abl4, \op-T0-cpy/iny ;
wire a1, dpc32_PCHADH, \A+B5 , ab12, net1238, \op-T2-branch , net1240, AxB7, adl2, \op-T+-ora/and/eor/adc ;
wire net1244, net1245, \op-shift-right , net1247, alua1, net1249, abl3, net1251, net1252, net1253;
wire net1254, net1255, net1256, net1257, net1258, \op-T4-ind-x , net1260, net1262, dpc2_XSB, net1264;
wire net1265, notdor5, net1267, \~DBZ , net1269, net1270, net1271, \notRdy0.phi1 , \op-T0 , net1274;
wire net1275, net1276, net1277, net1278, net1279, net1280, net1281, adl1, pipeUNK12, notidl3;
wire C01, net1286, sb2, notdor2, net1289, net1290, net1291, \op-T0-cli/sei , net1293, \PD-1xx000x0 ;
wire net1295, net1296, nmi, net1298, adl7, net1300, pchp5, idb3, net1303, net1304;
wire net1305, idl4, \~ABL6 , notaluvout, net1309, net1310, \op-T4-rti , net1312, \A+B3 , C67;
wire net1315, net1316, \~A.B7 , net1319, notir7, pipeUNK26, net1322, net1323, \op-T+-shift-a , net1325;
wire \~pclp5 , \~C78 , ir7, ir5, net1330, dpc26_ACDB, alua2, net1333, dpc35_PCHC, net1335;
wire sb6, \op-T0-cpx/cpy/inx/iny , net1338, net1339, ab2, net1341, \op-T0-acc , net1343, net1344, net1345;
wire net1346, net1347, net1348, db7, INTG, net1351, \~WR , net1353, net1354, \op-T0-cmp ;
wire net1356, net1357, net1358, pcl3, net1360, net1362, net1364, net1365, net1366, net1367;
wire net1368, net1369, Pout7, net1371, DC34, pipeT4out, NMIL, net1375, net1376, net1377;
wire net1378, net1379, net1380, \op-T3-jmp , \brk-done , net1383, ir2, \op-T5-mem-ind-idx , net1386, net1387;
wire net1388, net1389, net1390, net1391, net1392, db4, notir5, net1395, \op-T0-shift-a , net1397;
wire \~(A+B)7 , net1399, net1400, net1401, net1402, s0, net1404, dasb4, net1406, net1407;
wire net1408, net1409, \pd7.clearIR , net1411, net1412, net1413, alu3, dor6, net1416, net1417;
wire notdor6, \op-T0-cld/sed , \op-T0-lda , Pout2, net1422, net1423, net1424, \~C34 , net1426, net1427;
wire \op-T3-ind-x , abh0, \x-op-T3-plp/pla , \pipe~VEC , alub1, net1433, notx1, s7, pipeUNK03, adl4;
wire pipeUNK41, noty6, net1440, net1441, pipeUNK13, ab10, Pout1, net1445, net1446, net1447;
wire net1448, net1449, net1450, net1451, net1452, dor5, net1454, net1455, net1456, net1457;
wire pclp6, \~(AxB)6 , \pd6.clearIR , net1462, net1463, net1464, VEC0, \op-rol/ror , net1467, dpc5_SADL;
wire \~(AxB)5 , net1470, net1471, net1472, idb2, net1474, dasb3, \x-op-T0-bit , net1477, \op-T0-brk/rti ;
wire net1479, net1480, VEC1, \op-T+-iny/dey , net1483, noty2, notidl2, net1486, \op-T3-plp/pla , net1488;
wire net1489, notalu4, net1491, net1492, ab7, dasb7, net1495, pchp2, net1497, net1498;
wire net1499, net1500, net1501, abl2, idb5, \op-T0-and , net1505, \~C01 , net1507, net1508;
wire net1509, net1510, net1511, \op-T2-abs-y , \~ABL5 , net1514, net1515, notidl4, net1517, net1518;
wire net1519, \op-plp/pla , notx3, alua7, net1523, \op-T2-ind , \~(AxB)0 , net1526, net1527, net1528;
wire net1529, pipeUNK01, net1531, s3, net1533, net1534, alub7, clock1, notidl6, net1538;
wire adh7, \op-from-x , net1541, net1542, \x-op-T0-txa , BRtaken, net1545, net1546, net1547, net1548;
wire net1549, net1550, pch6, net1552, p2, net1554, net1555, net1556, \op-brk/rti , net1558;
wire net1559, net1560, notx7, \op-xy , net1563, \dpc41_DL/ADL , net1565, net1566, t3, net1568;
wire \x-op-T4-rti , net1570, \~C45 , net1572, net1573, net1574, net1575, ir3, pipeUNK15, net1578;
wire net1579, net1580, net1581, \op-T2-stack , net1583, net1584, net1585, net1586, \pd3.clearIR , net1588;
wire \op-T4-jmp , net1590, db6, net1592, net1593, net1594, net1595, net1596, idl0, net1598;
wire net1599, net1600, \op-sty/cpy-mem , net1602, nots4, net1604, net1605, net1606, pipeUNK14, net1608;
wire net1609, net1610, pcl7, \op-T4-rts , net1613, net1614, net1615, net1616, net1617, net1618;
wire net1619, net1620, net1621, \pd0.clearIR , \op-T0-eor , net1624, net1625, ir1, alua6, \~A.B0 ;
wire net1629, adl5, net1631, \~(A+B)5 , net1633, dor2, net1635, net1636, alu2, net1638;
wire net1639, noty7, net1641, net1642, net1643, net1644, alub4, \op-T+-bit , pclp7, x3;
wire net1649, net1650, adh2, pipeUNK30, a7, net1654, net1655, net1656, net1657, \op-T0-cpx/inx ;
wire net1659, net1660, net1661, net1662, \op-T+-inx , \op-T+-asl/rol-a , dpc16_EORS, net1667, net1668, pd6;
wire pch0, \pd2.clearIR , so, net1673, net1674, net1675, net1676, net1677, alub5, net1679;
wire alua3, net1681, net1682, net1683, net1684, net1685, net1686, net1687, net1688, \op-EORS ;
wire pd7, \~(A+B)2 , net1692, net1693, net1694, net1695, net1696, net1697, dpc24_ACSB, net1699;
wire dpc4_SSB, s4, net1703, dpc34_PCLC, net1705, net1706, net1707, \~op-T3-branch , net1709, \op-T+-cpx/cpy-imm/zp ;
wire net1711, net1712, pipeUNK35, net1714, net1715, net1716, net1717, net1718, net1719, net1720;
wire \op-branch-done , pchp0, net1723, net1724;

PULLUP pullup0 (.y(\op-T5-rts ));
PULLUP pullup3 (.y(net3));
PULLUP pullup4 (.y(\op-T0-tay ));
PULLUP pullup5 (.y(net5));
PULLUP pullup6 (.y(net6));
PULLUP pullup8 (.y(net8));
PULLUP pullup10 (.y(net10));
PULLUP pullup11 (.y(net11));
PULLUP pullup14 (.y(net14));
PULLUP pullup16 (.y(net16));
PULLUP pullup17 (.y(net17));
PULLUP pullup19 (.y(net19));
PULLUP pullup20 (.y(net20));
PULLUP pullup21 (.y(net21));
PULLUP pullup22 (.y(\~(AxBxC)2 ));
PULLUP pullup23 (.y(net23));
PULLUP pullup25 (.y(net25));
PULLUP pullup26 (.y(notir4));
PULLUP pullup27 (.y(pchp4));
PULLUP pullup29 (.y(net29));
PULLUP pullup31 (.y(net31));
PULLUP pullup33 (.y(\~pchp5 ));
PULLUP pullup34 (.y(net34));
PULLUP pullup35 (.y(net35));
PULLUP pullup36 (.y(net36));
PULLUP pullup38 (.y(net38));
PULLUP pullup39 (.y(\~pclp4 ));
PULLUP pullup46 (.y(net46));
PULLUP pullup53 (.y(\op-lsr/ror/dec/inc ));
PULLUP pullup58 (.y(\op-T3-abs-idx ));
PULLUP pullup60 (.y(\op-T3-ind-y ));
PULLUP pullup61 (.y(net61));
PULLUP pullup62 (.y(net62));
PULLUP pullup63 (.y(dor7));
PULLUP pullup65 (.y(\(AxB)4.~C34 ));
PULLUP pullup67 (.y(RESP));
PULLUP pullup70 (.y(net70));
PULLUP pullup71 (.y(net71));
PULLUP pullup72 (.y(pclp5));
PULLUP pullup75 (.y(net75));
PULLUP pullup76 (.y(\op-T0-dex ));
PULLUP pullup77 (.y(Pout6));
PULLUP pullup78 (.y(C34));
PULLUP pullup79 (.y(net79));
PULLUP pullup80 (.y(net80));
PULLUP pullup83 (.y(net83));
PULLUP pullup84 (.y(\op-T2-ind-x ));
PULLUP pullup89 (.y(rdy));
PULLUP pullup90 (.y(net90));
PULLUP pullup91 (.y(net91));
PULLUP pullup93 (.y(net93));
PULLUP pullup97 (.y(dor0));
PULLUP pullup104 (.y(net104));
PULLUP pullup105 (.y(net105));
PULLUP pullup108 (.y(net108));
PULLUP pullup109 (.y(net109));
PULLUP pullup110 (.y(\A+B2 ));
PULLUP pullup111 (.y(net111));
PULLUP pullup113 (.y(\~pchp1 ));
PULLUP pullup117 (.y(\A+B7 ));
PULLUP pullup118 (.y(net118));
PULLUP pullup120 (.y(\op-T3 ));
PULLUP pullup122 (.y(net122));
PULLUP pullup123 (.y(net123));
PULLUP pullup124 (.y(\~pchp3 ));
PULLUP pullup125 (.y(\PD-n-0xx0xx0x ));
PULLUP pullup127 (.y(net127));
PULLUP pullup128 (.y(net128));
PULLUP pullup130 (.y(net130));
PULLUP pullup131 (.y(\op-T0-pla ));
PULLUP pullup132 (.y(net132));
PULLUP pullup133 (.y(net133));
PULLUP pullup134 (.y(net134));
PULLUP pullup139 (.y(net139));
PULLUP pullup141 (.y(pchp3));
PULLUP pullup142 (.y(C45));
PULLUP pullup143 (.y(\~(A+B)0 ));
PULLUP pullup145 (.y(\op-sta/cmp ));
PULLUP pullup146 (.y(net146));
PULLUP pullup149 (.y(net149));
PULLUP pullup152 (.y(net152));
PULLUP pullup154 (.y(net154));
PULLUP pullup155 (.y(\~(A+B)1 ));
PULLUP pullup156 (.y(clock2));
PULLUP pullup157 (.y(\op-T2-stack-access ));
PULLUP pullup160 (.y(net160));
PULLUP pullup161 (.y(net161));
PULLUP pullup163 (.y(net163));
PULLUP pullup167 (.y(\op-T0-tax ));
PULLUP pullup168 (.y(net168));
PULLUP pullup169 (.y(net169));
PULLUP pullup172 (.y(net172));
PULLUP pullup174 (.y(\(AxB)6.~C56 ));
PULLUP pullup176 (.y(net176));
PULLUP pullup177 (.y(\~(AxB)7 ));
PULLUP pullup178 (.y(abl6));
PULLUP pullup179 (.y(\op-T0-txa ));
PULLUP pullup180 (.y(net180));
PULLUP pullup182 (.y(net182));
PULLUP pullup184 (.y(noty3));
PULLUP pullup187 (.y(notRnWprepad));
PULLUP pullup188 (.y(net188));
PULLUP pullup191 (.y(net191));
PULLUP pullup192 (.y(net192));
PULLUP pullup193 (.y(\(AxB)2.~C12 ));
PULLUP pullup194 (.y(notir0));
PULLUP pullup196 (.y(net196));
PULLUP pullup198 (.y(net198));
PULLUP pullup200 (.y(net200));
PULLUP pullup201 (.y(net201));
PULLUP pullup204 (.y(\op-T2-ADL/ADD ));
PULLUP pullup206 (.y(\~alucout ));
PULLUP pullup207 (.y(net207));
PULLUP pullup208 (.y(pclp4));
PULLUP pullup209 (.y(pchp1));
PULLUP pullup212 (.y(net212));
PULLUP pullup213 (.y(net213));
PULLUP pullup216 (.y(\DA-AB2 ));
PULLUP pullup217 (.y(\0/ADL0 ));
PULLUP pullup218 (.y(net218));
PULLUP pullup219 (.y(\op-T2-mem-zp ));
PULLUP pullup220 (.y(net220));
PULLUP pullup221 (.y(net221));
PULLUP pullup224 (.y(net224));
PULLUP pullup225 (.y(net225));
PULLUP pullup227 (.y(net227));
PULLUP pullup228 (.y(net228));
PULLUP pullup229 (.y(dpc28_0ADH0));
PULLUP pullup231 (.y(net231));
PULLUP pullup232 (.y(net232));
PULLUP pullup233 (.y(net233));
PULLUP pullup234 (.y(abl5));
PULLUP pullup236 (.y(net236));
PULLUP pullup238 (.y(net238));
PULLUP pullup240 (.y(idl5));
PULLUP pullup241 (.y(net241));
PULLUP pullup242 (.y(net242));
PULLUP pullup243 (.y(net243));
PULLUP pullup244 (.y(\op-ror ));
PULLUP pullup245 (.y(\op-T0-txs ));
PULLUP pullup249 (.y(net249));
PULLUP pullup251 (.y(net251));
PULLUP pullup252 (.y(\~op-set-C ));
PULLUP pullup253 (.y(net253));
PULLUP pullup254 (.y(net254));
PULLUP pullup255 (.y(net255));
PULLUP pullup256 (.y(net256));
PULLUP pullup257 (.y(\op-T0-tya ));
PULLUP pullup258 (.y(\op-T2-idx-x-xy ));
PULLUP pullup259 (.y(\op-jsr ));
PULLUP pullup260 (.y(net260));
PULLUP pullup261 (.y(net261));
PULLUP pullup262 (.y(net262));
PULLUP pullup263 (.y(dasb5));
PULLUP pullup264 (.y(\~NMIG ));
PULLUP pullup267 (.y(net267));
PULLUP pullup269 (.y(net269));
PULLUP pullup270 (.y(net270));
PULLUP pullup271 (.y(\op-T0-jsr ));
PULLUP pullup272 (.y(net272));
PULLUP pullup273 (.y(\op-T2-abs-access ));
PULLUP pullup274 (.y(\~(AxBxC)3 ));
PULLUP pullup275 (.y(net275));
PULLUP pullup278 (.y(net278));
PULLUP pullup279 (.y(net279));
PULLUP pullup280 (.y(net280));
PULLUP pullup281 (.y(\op-T4-mem-abs-idx ));
PULLUP pullup282 (.y(net282));
PULLUP pullup284 (.y(net284));
PULLUP pullup285 (.y(\op-T2-zp/zp-idx ));
PULLUP pullup286 (.y(\op-T0-tay/ldy-not-idx ));
PULLUP pullup287 (.y(abh2));
PULLUP pullup288 (.y(net288));
PULLUP pullup291 (.y(net291));
PULLUP pullup293 (.y(net293));
PULLUP pullup295 (.y(\~(AxB1).C01 ));
PULLUP pullup297 (.y(\~NMIP ));
PULLUP pullup299 (.y(net299));
PULLUP pullup300 (.y(net300));
PULLUP pullup301 (.y(\op-T+-cmp ));
PULLUP pullup302 (.y(\PD-xxx010x1 ));
PULLUP pullup303 (.y(\op-T0-bit ));
PULLUP pullup306 (.y(net306));
PULLUP pullup307 (.y(net307));
PULLUP pullup308 (.y(\~(AxB)4 ));
PULLUP pullup309 (.y(\op-T2-jmp-abs ));
PULLUP pullup311 (.y(net311));
PULLUP pullup312 (.y(net312));
PULLUP pullup314 (.y(alu5));
PULLUP pullup317 (.y(net317));
PULLUP pullup318 (.y(net318));
PULLUP pullup319 (.y(net319));
PULLUP pullup320 (.y(net320));
PULLUP pullup321 (.y(net321));
PULLUP pullup324 (.y(\op-inc/nop ));
PULLUP pullup326 (.y(net326));
PULLUP pullup327 (.y(net327));
PULLUP pullup328 (.y(ir0));
PULLUP pullup329 (.y(net329));
PULLUP pullup330 (.y(net330));
PULLUP pullup331 (.y(alu6));
PULLUP pullup332 (.y(net332));
PULLUP pullup333 (.y(DC78));
PULLUP pullup334 (.y(net334));
PULLUP pullup335 (.y(net335));
PULLUP pullup336 (.y(\~A.B6 ));
PULLUP pullup337 (.y(ir6));
PULLUP pullup340 (.y(net340));
PULLUP pullup341 (.y(\op-T4 ));
PULLUP pullup342 (.y(\x-op-T3-ind-y ));
PULLUP pullup344 (.y(net344));
PULLUP pullup345 (.y(net345));
PULLUP pullup347 (.y(net347));
PULLUP pullup350 (.y(\~A.B3 ));
PULLUP pullup351 (.y(net351));
PULLUP pullup352 (.y(\op-T4-brk ));
PULLUP pullup354 (.y(\op-T4-abs-idx ));
PULLUP pullup355 (.y(net355));
PULLUP pullup358 (.y(net358));
PULLUP pullup365 (.y(\PD-0xx0xx0x ));
PULLUP pullup366 (.y(net366));
PULLUP pullup368 (.y(net368));
PULLUP pullup370 (.y(\op-T5-brk ));
PULLUP pullup371 (.y(\~(AxBxC)0 ));
PULLUP pullup372 (.y(net372));
PULLUP pullup374 (.y(net374));
PULLUP pullup376 (.y(abl1));
PULLUP pullup378 (.y(net378));
PULLUP pullup379 (.y(\dpc36_~IPC ));
PULLUP pullup382 (.y(\op-T0-iny/dey ));
PULLUP pullup383 (.y(net383));
PULLUP pullup384 (.y(net384));
PULLUP pullup385 (.y(net385));
PULLUP pullup386 (.y(net386));
PULLUP pullup388 (.y(net388));
PULLUP pullup389 (.y(net389));
PULLUP pullup390 (.y(net390));
PULLUP pullup391 (.y(idl7));
PULLUP pullup392 (.y(net392));
PULLUP pullup396 (.y(net396));
PULLUP pullup397 (.y(net397));
PULLUP pullup400 (.y(net400));
PULLUP pullup401 (.y(alu0));
PULLUP pullup403 (.y(\op-T0-ora ));
PULLUP pullup404 (.y(\~(A+B)4 ));
PULLUP pullup409 (.y(net409));
PULLUP pullup410 (.y(net410));
PULLUP pullup412 (.y(notalucout));
PULLUP pullup419 (.y(net419));
PULLUP pullup420 (.y(net420));
PULLUP pullup422 (.y(abh3));
PULLUP pullup423 (.y(net423));
PULLUP pullup424 (.y(net424));
PULLUP pullup425 (.y(AxB1));
PULLUP pullup427 (.y(\~C56 ));
PULLUP pullup428 (.y(net428));
PULLUP pullup432 (.y(net432));
PULLUP pullup434 (.y(\op-rmw ));
PULLUP pullup436 (.y(net436));
PULLUP pullup439 (.y(Pout3));
PULLUP pullup440 (.y(net440));
PULLUP pullup441 (.y(net441));
PULLUP pullup442 (.y(net442));
PULLUP pullup444 (.y(dor3));
PULLUP pullup445 (.y(net445));
PULLUP pullup446 (.y(\op-T5-rti/rts ));
PULLUP pullup447 (.y(\x-op-T3-abs-idx ));
PULLUP pullup450 (.y(dasb2));
PULLUP pullup453 (.y(net453));
PULLUP pullup457 (.y(net457));
PULLUP pullup458 (.y(net458));
PULLUP pullup461 (.y(\x-op-T4-ind-y ));
PULLUP pullup462 (.y(net462));
PULLUP pullup464 (.y(idl3));
PULLUP pullup465 (.y(\~~alucout ));
PULLUP pullup466 (.y(net466));
PULLUP pullup467 (.y(net467));
PULLUP pullup468 (.y(net468));
PULLUP pullup470 (.y(net470));
PULLUP pullup472 (.y(net472));
PULLUP pullup473 (.y(net473));
PULLUP pullup474 (.y(net474));
PULLUP pullup476 (.y(net476));
PULLUP pullup477 (.y(\~A.B5 ));
PULLUP pullup478 (.y(net478));
PULLUP pullup479 (.y(net479));
PULLUP pullup480 (.y(net480));
PULLUP pullup481 (.y(pclp2));
PULLUP pullup484 (.y(net484));
PULLUP pullup485 (.y(notx4));
PULLUP pullup486 (.y(\~(AxBxC)5 ));
PULLUP pullup487 (.y(\op-T2-brk ));
PULLUP pullup488 (.y(pclp0));
PULLUP pullup489 (.y(abh7));
PULLUP pullup490 (.y(net490));
PULLUP pullup491 (.y(net491));
PULLUP pullup492 (.y(\op-T4-ind-y ));
PULLUP pullup494 (.y(net494));
PULLUP pullup496 (.y(net496));
PULLUP pullup499 (.y(net499));
PULLUP pullup500 (.y(C56));
PULLUP pullup501 (.y(net501));
PULLUP pullup503 (.y(net503));
PULLUP pullup504 (.y(net504));
PULLUP pullup505 (.y(C12));
PULLUP pullup506 (.y(net506));
PULLUP pullup507 (.y(net507));
PULLUP pullup510 (.y(net510));
PULLUP pullup513 (.y(net513));
PULLUP pullup515 (.y(net515));
PULLUP pullup516 (.y(\DA-AxB2 ));
PULLUP pullup517 (.y(\op-store ));
PULLUP pullup518 (.y(net518));
PULLUP pullup519 (.y(net519));
PULLUP pullup522 (.y(\op-ORS ));
PULLUP pullup523 (.y(net523));
PULLUP pullup525 (.y(net525));
PULLUP pullup528 (.y(\xx-op-T5-jsr ));
PULLUP pullup531 (.y(net531));
PULLUP pullup532 (.y(\~(AxBxC)7 ));
PULLUP pullup533 (.y(net533));
PULLUP pullup535 (.y(\~pchp7 ));
PULLUP pullup538 (.y(net538));
PULLUP pullup540 (.y(\pd4.clearIR ));
PULLUP pullup543 (.y(net543));
PULLUP pullup544 (.y(net544));
PULLUP pullup546 (.y(\op-shift ));
PULLUP pullup548 (.y(net548));
PULLUP pullup550 (.y(net550));
PULLUP pullup551 (.y(net551));
PULLUP pullup552 (.y(\op-T0-php/pha ));
PULLUP pullup553 (.y(net553));
PULLUP pullup555 (.y(\(AxB)0.~C0in ));
PULLUP pullup556 (.y(net556));
PULLUP pullup564 (.y(net564));
PULLUP pullup565 (.y(noty4));
PULLUP pullup566 (.y(net566));
PULLUP pullup567 (.y(abl7));
PULLUP pullup568 (.y(net568));
PULLUP pullup570 (.y(net570));
PULLUP pullup571 (.y(net571));
PULLUP pullup572 (.y(net572));
PULLUP pullup575 (.y(\op-T0-adc/sbc ));
PULLUP pullup578 (.y(net578));
PULLUP pullup579 (.y(\op-T3-jsr ));
PULLUP pullup582 (.y(net582));
PULLUP pullup583 (.y(net583));
PULLUP pullup586 (.y(net586));
PULLUP pullup587 (.y(net587));
PULLUP pullup588 (.y(net588));
PULLUP pullup592 (.y(\~C67 ));
PULLUP pullup593 (.y(net593));
PULLUP pullup594 (.y(\op-T0-jmp ));
PULLUP pullup595 (.y(net595));
PULLUP pullup600 (.y(net600));
PULLUP pullup602 (.y(net602));
PULLUP pullup603 (.y(net603));
PULLUP pullup604 (.y(net604));
PULLUP pullup606 (.y(alu4));
PULLUP pullup607 (.y(\op-T3-mem-abs ));
PULLUP pullup608 (.y(net608));
PULLUP pullup609 (.y(net609));
PULLUP pullup611 (.y(net611));
PULLUP pullup613 (.y(net613));
PULLUP pullup616 (.y(net616));
PULLUP pullup617 (.y(net617));
PULLUP pullup618 (.y(net618));
PULLUP pullup620 (.y(net620));
PULLUP pullup623 (.y(\DA-C01 ));
PULLUP pullup624 (.y(net624));
PULLUP pullup625 (.y(net625));
PULLUP pullup626 (.y(\branch-back ));
PULLUP pullup628 (.y(net628));
PULLUP pullup629 (.y(net629));
PULLUP pullup630 (.y(net630));
PULLUP pullup631 (.y(net631));
PULLUP pullup632 (.y(net632));
PULLUP pullup636 (.y(net636));
PULLUP pullup637 (.y(net637));
PULLUP pullup638 (.y(net638));
PULLUP pullup640 (.y(AxB3));
PULLUP pullup641 (.y(net641));
PULLUP pullup645 (.y(net645));
PULLUP pullup646 (.y(net646));
PULLUP pullup647 (.y(net647));
PULLUP pullup649 (.y(\~(A+B)3 ));
PULLUP pullup651 (.y(\~(AxBxC)4 ));
PULLUP pullup652 (.y(pchp6));
PULLUP pullup658 (.y(net658));
PULLUP pullup660 (.y(\op-T3-branch ));
PULLUP pullup662 (.y(net662));
PULLUP pullup664 (.y(net664));
PULLUP pullup665 (.y(\op-T0-ldy-mem ));
PULLUP pullup667 (.y(\pd5.clearIR ));
PULLUP pullup669 (.y(net669));
PULLUP pullup670 (.y(net670));
PULLUP pullup673 (.y(net673));
PULLUP pullup674 (.y(net674));
PULLUP pullup677 (.y(\op-T3-abs/idx/ind ));
PULLUP pullup678 (.y(net678));
PULLUP pullup679 (.y(dasb6));
PULLUP pullup681 (.y(\~A.B2 ));
PULLUP pullup682 (.y(\op-T0-tsx ));
PULLUP pullup686 (.y(\0/ADL1 ));
PULLUP pullup687 (.y(Pout0));
PULLUP pullup689 (.y(net689));
PULLUP pullup690 (.y(t4));
PULLUP pullup691 (.y(\op-asl/rol ));
PULLUP pullup692 (.y(net692));
PULLUP pullup693 (.y(\A+B0 ));
PULLUP pullup694 (.y(net694));
PULLUP pullup695 (.y(net695));
PULLUP pullup696 (.y(net696));
PULLUP pullup699 (.y(\~DA-ADD2 ));
PULLUP pullup700 (.y(net700));
PULLUP pullup701 (.y(\~(AxB)2 ));
PULLUP pullup702 (.y(notir1));
PULLUP pullup708 (.y(net708));
PULLUP pullup709 (.y(net709));
PULLUP pullup712 (.y(\op-T2-jsr ));
PULLUP pullup713 (.y(abh1));
PULLUP pullup714 (.y(net714));
PULLUP pullup715 (.y(net715));
PULLUP pullup717 (.y(net717));
PULLUP pullup718 (.y(net718));
PULLUP pullup720 (.y(net720));
PULLUP pullup721 (.y(net721));
PULLUP pullup723 (.y(pclp3));
PULLUP pullup725 (.y(\dpc22_~DSA ));
PULLUP pullup726 (.y(net726));
PULLUP pullup728 (.y(net728));
PULLUP pullup730 (.y(notx6));
PULLUP pullup731 (.y(\~pclp6 ));
PULLUP pullup732 (.y(net732));
PULLUP pullup733 (.y(net733));
PULLUP pullup735 (.y(net735));
PULLUP pullup739 (.y(net739));
PULLUP pullup743 (.y(net743));
PULLUP pullup744 (.y(DBZ));
PULLUP pullup746 (.y(dor1));
PULLUP pullup747 (.y(net747));
PULLUP pullup748 (.y(net748));
PULLUP pullup750 (.y(\op-T2-php ));
PULLUP pullup753 (.y(net753));
PULLUP pullup754 (.y(net754));
PULLUP pullup755 (.y(net755));
PULLUP pullup757 (.y(net757));
PULLUP pullup761 (.y(net761));
PULLUP pullup762 (.y(net762));
PULLUP pullup763 (.y(net763));
PULLUP pullup764 (.y(\op-jmp ));
PULLUP pullup765 (.y(alu7));
PULLUP pullup767 (.y(net767));
PULLUP pullup769 (.y(net769));
PULLUP pullup770 (.y(\notRdy0.delay ));
PULLUP pullup771 (.y(\branch-back.phi1 ));
PULLUP pullup772 (.y(net772));
PULLUP pullup773 (.y(net773));
PULLUP pullup774 (.y(net774));
PULLUP pullup775 (.y(abh5));
PULLUP pullup776 (.y(\op-T5-jsr ));
PULLUP pullup778 (.y(ONEBYTE));
PULLUP pullup779 (.y(net779));
PULLUP pullup781 (.y(net781));
PULLUP pullup782 (.y(net782));
PULLUP pullup783 (.y(net783));
PULLUP pullup784 (.y(\op-T5-rti ));
PULLUP pullup786 (.y(\op-T+-dex ));
PULLUP pullup787 (.y(\op-T0-sbc ));
PULLUP pullup788 (.y(\op-T2 ));
PULLUP pullup789 (.y(net789));
PULLUP pullup790 (.y(net790));
PULLUP pullup791 (.y(\op-push/pull ));
PULLUP pullup795 (.y(net795));
PULLUP pullup797 (.y(net797));
PULLUP pullup800 (.y(net800));
PULLUP pullup803 (.y(\A+B6 ));
PULLUP pullup804 (.y(\op-T4-brk/jsr ));
PULLUP pullup807 (.y(net807));
PULLUP pullup808 (.y(alurawcout));
PULLUP pullup809 (.y(\pd1.clearIR ));
PULLUP pullup810 (.y(net810));
PULLUP pullup811 (.y(net811));
PULLUP pullup812 (.y(net812));
PULLUP pullup813 (.y(net813));
PULLUP pullup815 (.y(net815));
PULLUP pullup817 (.y(\~(AxB5).C45 ));
PULLUP pullup818 (.y(net818));
PULLUP pullup819 (.y(net819));
PULLUP pullup822 (.y(\op-T+-adc/sbc ));
PULLUP pullup824 (.y(net824));
PULLUP pullup827 (.y(D1x1));
PULLUP pullup830 (.y(net830));
PULLUP pullup831 (.y(net831));
PULLUP pullup834 (.y(net834));
PULLUP pullup837 (.y(net837));
PULLUP pullup838 (.y(net838));
PULLUP pullup839 (.y(net839));
PULLUP pullup840 (.y(\~op-branch-bit6 ));
PULLUP pullup841 (.y(\~A.B1 ));
PULLUP pullup842 (.y(net842));
PULLUP pullup844 (.y(net844));
PULLUP pullup845 (.y(net845));
PULLUP pullup846 (.y(net846));
PULLUP pullup847 (.y(net847));
PULLUP pullup849 (.y(net849));
PULLUP pullup850 (.y(net850));
PULLUP pullup851 (.y(\~TWOCYCLE ));
PULLUP pullup852 (.y(net852));
PULLUP pullup853 (.y(net853));
PULLUP pullup854 (.y(net854));
PULLUP pullup857 (.y(\op-rti/rts ));
PULLUP pullup860 (.y(\~(AxB3).C23 ));
PULLUP pullup861 (.y(net861));
PULLUP pullup862 (.y(net862));
PULLUP pullup867 (.y(net867));
PULLUP pullup870 (.y(idl1));
PULLUP pullup871 (.y(net871));
PULLUP pullup872 (.y(alu1));
PULLUP pullup875 (.y(net875));
PULLUP pullup876 (.y(net876));
PULLUP pullup877 (.y(net877));
PULLUP pullup879 (.y(fetch));
PULLUP pullup880 (.y(net880));
PULLUP pullup882 (.y(net882));
PULLUP pullup883 (.y(net883));
PULLUP pullup884 (.y(\~(AxB)3 ));
PULLUP pullup885 (.y(net885));
PULLUP pullup888 (.y(\~IRQP ));
PULLUP pullup889 (.y(net889));
PULLUP pullup890 (.y(notx2));
PULLUP pullup895 (.y(notir6));
PULLUP pullup896 (.y(net896));
PULLUP pullup901 (.y(\~DA-ADD1 ));
PULLUP pullup904 (.y(\op-T3-mem-zp-idx ));
PULLUP pullup905 (.y(net905));
PULLUP pullup906 (.y(net906));
PULLUP pullup909 (.y(t5));
PULLUP pullup910 (.y(alucin));
PULLUP pullup913 (.y(net913));
PULLUP pullup916 (.y(net916));
PULLUP pullup917 (.y(net917));
PULLUP pullup918 (.y(\A+B4 ));
PULLUP pullup919 (.y(net919));
PULLUP pullup920 (.y(net920));
PULLUP pullup923 (.y(net923));
PULLUP pullup925 (.y(\~op-store ));
PULLUP pullup926 (.y(RESG));
PULLUP pullup928 (.y(net928));
PULLUP pullup929 (.y(net929));
PULLUP pullup930 (.y(net930));
PULLUP pullup931 (.y(net931));
PULLUP pullup932 (.y(\op-T2-php/pha ));
PULLUP pullup933 (.y(net933));
PULLUP pullup934 (.y(\op-SRS ));
PULLUP pullup935 (.y(net935));
PULLUP pullup936 (.y(net936));
PULLUP pullup937 (.y(net937));
PULLUP pullup938 (.y(aluvout));
PULLUP pullup944 (.y(net944));
PULLUP pullup946 (.y(net946));
PULLUP pullup947 (.y(net947));
PULLUP pullup950 (.y(\op-T+-cpx/cpy-abs ));
PULLUP pullup951 (.y(net951));
PULLUP pullup952 (.y(net952));
PULLUP pullup953 (.y(\~(AxB)1 ));
PULLUP pullup954 (.y(net954));
PULLUP pullup956 (.y(net956));
PULLUP pullup958 (.y(net958));
PULLUP pullup959 (.y(net959));
PULLUP pullup961 (.y(net961));
PULLUP pullup962 (.y(net962));
PULLUP pullup964 (.y(net964));
PULLUP pullup965 (.y(\~(AxBxC)1 ));
PULLUP pullup966 (.y(net966));
PULLUP pullup967 (.y(nnT2BR));
PULLUP pullup969 (.y(net969));
PULLUP pullup971 (.y(t2));
PULLUP pullup973 (.y(net973));
PULLUP pullup975 (.y(net975));
PULLUP pullup976 (.y(pclp1));
PULLUP pullup979 (.y(net979));
PULLUP pullup980 (.y(net980));
PULLUP pullup981 (.y(noty5));
PULLUP pullup983 (.y(net983));
PULLUP pullup985 (.y(\op-T0-ldx/tax/tsx ));
PULLUP pullup986 (.y(net986));
PULLUP pullup987 (.y(notx0));
PULLUP pullup988 (.y(net988));
PULLUP pullup990 (.y(net990));
PULLUP pullup992 (.y(net992));
PULLUP pullup995 (.y(net995));
PULLUP pullup996 (.y(irline3));
PULLUP pullup997 (.y(abh6));
PULLUP pullup998 (.y(net998));
PULLUP pullup1002 (.y(net1002));
PULLUP pullup1003 (.y(\~C23 ));
PULLUP pullup1006 (.y(\op-implied ));
PULLUP pullup1007 (.y(net1007));
PULLUP pullup1009 (.y(dasb1));
PULLUP pullup1010 (.y(net1010));
PULLUP pullup1016 (.y(net1016));
PULLUP pullup1017 (.y(notx5));
PULLUP pullup1018 (.y(net1018));
PULLUP pullup1019 (.y(\PD-xxxx10x0 ));
PULLUP pullup1021 (.y(\A+B1 ));
PULLUP pullup1023 (.y(C23));
PULLUP pullup1024 (.y(net1024));
PULLUP pullup1025 (.y(noty0));
PULLUP pullup1026 (.y(net1026));
PULLUP pullup1028 (.y(net1028));
PULLUP pullup1031 (.y(\op-T3-stack/bit/jmp ));
PULLUP pullup1032 (.y(NMIP));
PULLUP pullup1033 (.y(net1033));
PULLUP pullup1034 (.y(net1034));
PULLUP pullup1035 (.y(\~DBE ));
PULLUP pullup1037 (.y(net1037));
PULLUP pullup1038 (.y(net1038));
PULLUP pullup1039 (.y(net1039));
PULLUP pullup1042 (.y(H1x1));
PULLUP pullup1043 (.y(net1043));
PULLUP pullup1044 (.y(net1044));
PULLUP pullup1045 (.y(net1045));
PULLUP pullup1046 (.y(net1046));
PULLUP pullup1047 (.y(net1047));
PULLUP pullup1048 (.y(\~op-branch-done ));
PULLUP pullup1050 (.y(\x-op-push/pull ));
PULLUP pullup1052 (.y(\x-op-jmp ));
PULLUP pullup1054 (.y(net1054));
PULLUP pullup1055 (.y(net1055));
PULLUP pullup1056 (.y(net1056));
PULLUP pullup1057 (.y(\op-T2-abs ));
PULLUP pullup1063 (.y(\~A.B4 ));
PULLUP pullup1065 (.y(net1065));
PULLUP pullup1066 (.y(idl2));
PULLUP pullup1067 (.y(net1067));
PULLUP pullup1069 (.y(net1069));
PULLUP pullup1070 (.y(net1070));
PULLUP pullup1073 (.y(net1073));
PULLUP pullup1074 (.y(\op-T0-shift-right-a ));
PULLUP pullup1075 (.y(net1075));
PULLUP pullup1077 (.y(clearIR));
PULLUP pullup1079 (.y(\~pclp2 ));
PULLUP pullup1081 (.y(net1081));
PULLUP pullup1082 (.y(net1082));
PULLUP pullup1083 (.y(net1083));
PULLUP pullup1084 (.y(\~(A+B)6 ));
PULLUP pullup1085 (.y(net1085));
PULLUP pullup1086 (.y(\op-T2-pha ));
PULLUP pullup1087 (.y(net1087));
PULLUP pullup1088 (.y(dor4));
PULLUP pullup1089 (.y(net1089));
PULLUP pullup1090 (.y(net1090));
PULLUP pullup1091 (.y(net1091));
PULLUP pullup1093 (.y(net1093));
PULLUP pullup1094 (.y(net1094));
PULLUP pullup1096 (.y(abl0));
PULLUP pullup1097 (.y(net1097));
PULLUP pullup1099 (.y(net1099));
PULLUP pullup1101 (.y(net1101));
PULLUP pullup1106 (.y(net1106));
PULLUP pullup1107 (.y(net1107));
PULLUP pullup1109 (.y(net1109));
PULLUP pullup1110 (.y(\branch-forward.phi1 ));
PULLUP pullup1111 (.y(net1111));
PULLUP pullup1112 (.y(ir4));
PULLUP pullup1114 (.y(\op-T0-clc/sec ));
PULLUP pullup1115 (.y(net1115));
PULLUP pullup1116 (.y(idl6));
PULLUP pullup1117 (.y(net1117));
PULLUP pullup1119 (.y(Pout4));
PULLUP pullup1120 (.y(net1120));
PULLUP pullup1122 (.y(\~C12 ));
PULLUP pullup1125 (.y(notir3));
PULLUP pullup1129 (.y(net1129));
PULLUP pullup1130 (.y(net1130));
PULLUP pullup1133 (.y(net1133));
PULLUP pullup1134 (.y(\~VEC ));
PULLUP pullup1135 (.y(net1135));
PULLUP pullup1137 (.y(net1137));
PULLUP pullup1138 (.y(noty1));
PULLUP pullup1141 (.y(net1141));
PULLUP pullup1143 (.y(abh4));
PULLUP pullup1144 (.y(\DA-C45 ));
PULLUP pullup1145 (.y(net1145));
PULLUP pullup1146 (.y(alucout));
PULLUP pullup1153 (.y(net1153));
PULLUP pullup1154 (.y(net1154));
PULLUP pullup1155 (.y(\x-op-T+-adc/sbc ));
PULLUP pullup1157 (.y(net1157));
PULLUP pullup1159 (.y(net1159));
PULLUP pullup1164 (.y(\op-clv ));
PULLUP pullup1165 (.y(notalucin));
PULLUP pullup1166 (.y(net1166));
PULLUP pullup1168 (.y(\op-T5-ind-y ));
PULLUP pullup1169 (.y(net1169));
PULLUP pullup1170 (.y(net1170));
PULLUP pullup1173 (.y(\x-op-T0-tya ));
PULLUP pullup1174 (.y(\~op-branch-bit7 ));
PULLUP pullup1175 (.y(net1175));
PULLUP pullup1178 (.y(net1178));
PULLUP pullup1179 (.y(net1179));
PULLUP pullup1180 (.y(net1180));
PULLUP pullup1181 (.y(net1181));
PULLUP pullup1182 (.y(notir2));
PULLUP pullup1184 (.y(net1184));
PULLUP pullup1185 (.y(\short-circuit-idx-add ));
PULLUP pullup1187 (.y(net1187));
PULLUP pullup1190 (.y(net1190));
PULLUP pullup1192 (.y(net1192));
PULLUP pullup1193 (.y(\0/ADL2 ));
PULLUP pullup1194 (.y(net1194));
PULLUP pullup1195 (.y(net1195));
PULLUP pullup1196 (.y(\op-SUMS ));
PULLUP pullup1197 (.y(\~(AxBxC)6 ));
PULLUP pullup1199 (.y(net1199));
PULLUP pullup1200 (.y(DBNeg));
PULLUP pullup1202 (.y(net1202));
PULLUP pullup1204 (.y(\op-T2-ind-y ));
PULLUP pullup1205 (.y(net1205));
PULLUP pullup1206 (.y(pchp7));
PULLUP pullup1209 (.y(net1209));
PULLUP pullup1210 (.y(\op-T5-ind-x ));
PULLUP pullup1211 (.y(net1211));
PULLUP pullup1213 (.y(net1213));
PULLUP pullup1214 (.y(net1214));
PULLUP pullup1215 (.y(net1215));
PULLUP pullup1217 (.y(\~(AxB7).C67 ));
PULLUP pullup1218 (.y(net1218));
PULLUP pullup1219 (.y(net1219));
PULLUP pullup1220 (.y(AxB5));
PULLUP pullup1222 (.y(net1222));
PULLUP pullup1223 (.y(net1223));
PULLUP pullup1224 (.y(net1224));
PULLUP pullup1225 (.y(net1225));
PULLUP pullup1226 (.y(\op-T0-plp ));
PULLUP pullup1227 (.y(\~pclp0 ));
PULLUP pullup1228 (.y(\op-ANDS ));
PULLUP pullup1229 (.y(net1229));
PULLUP pullup1230 (.y(net1230));
PULLUP pullup1231 (.y(net1231));
PULLUP pullup1232 (.y(abl4));
PULLUP pullup1233 (.y(\op-T0-cpy/iny ));
PULLUP pullup1236 (.y(\A+B5 ));
PULLUP pullup1238 (.y(net1238));
PULLUP pullup1239 (.y(\op-T2-branch ));
PULLUP pullup1240 (.y(net1240));
PULLUP pullup1241 (.y(AxB7));
PULLUP pullup1243 (.y(\op-T+-ora/and/eor/adc ));
PULLUP pullup1244 (.y(net1244));
PULLUP pullup1245 (.y(net1245));
PULLUP pullup1246 (.y(\op-shift-right ));
PULLUP pullup1250 (.y(abl3));
PULLUP pullup1251 (.y(net1251));
PULLUP pullup1253 (.y(net1253));
PULLUP pullup1255 (.y(net1255));
PULLUP pullup1256 (.y(net1256));
PULLUP pullup1257 (.y(net1257));
PULLUP pullup1258 (.y(net1258));
PULLUP pullup1259 (.y(\op-T4-ind-x ));
PULLUP pullup1260 (.y(net1260));
PULLUP pullup1262 (.y(net1262));
PULLUP pullup1265 (.y(net1265));
PULLUP pullup1267 (.y(net1267));
PULLUP pullup1268 (.y(\~DBZ ));
PULLUP pullup1270 (.y(net1270));
PULLUP pullup1271 (.y(net1271));
PULLUP pullup1273 (.y(\op-T0 ));
PULLUP pullup1275 (.y(net1275));
PULLUP pullup1277 (.y(net1277));
PULLUP pullup1281 (.y(net1281));
PULLUP pullup1285 (.y(C01));
PULLUP pullup1286 (.y(net1286));
PULLUP pullup1289 (.y(net1289));
PULLUP pullup1290 (.y(net1290));
PULLUP pullup1292 (.y(\op-T0-cli/sei ));
PULLUP pullup1293 (.y(net1293));
PULLUP pullup1294 (.y(\PD-1xx000x0 ));
PULLUP pullup1295 (.y(net1295));
PULLUP pullup1301 (.y(pchp5));
PULLUP pullup1303 (.y(net1303));
PULLUP pullup1304 (.y(net1304));
PULLUP pullup1305 (.y(net1305));
PULLUP pullup1306 (.y(idl4));
PULLUP pullup1308 (.y(notaluvout));
PULLUP pullup1309 (.y(net1309));
PULLUP pullup1311 (.y(\op-T4-rti ));
PULLUP pullup1312 (.y(net1312));
PULLUP pullup1313 (.y(\A+B3 ));
PULLUP pullup1314 (.y(C67));
PULLUP pullup1315 (.y(net1315));
PULLUP pullup1316 (.y(net1316));
PULLUP pullup1318 (.y(\~A.B7 ));
PULLUP pullup1319 (.y(net1319));
PULLUP pullup1320 (.y(notir7));
PULLUP pullup1323 (.y(net1323));
PULLUP pullup1324 (.y(\op-T+-shift-a ));
PULLUP pullup1327 (.y(\~C78 ));
PULLUP pullup1328 (.y(ir7));
PULLUP pullup1329 (.y(ir5));
PULLUP pullup1334 (.y(dpc35_PCHC));
PULLUP pullup1335 (.y(net1335));
PULLUP pullup1337 (.y(\op-T0-cpx/cpy/inx/iny ));
PULLUP pullup1339 (.y(net1339));
PULLUP pullup1342 (.y(\op-T0-acc ));
PULLUP pullup1343 (.y(net1343));
PULLUP pullup1344 (.y(net1344));
PULLUP pullup1345 (.y(net1345));
PULLUP pullup1346 (.y(net1346));
PULLUP pullup1347 (.y(net1347));
PULLUP pullup1350 (.y(INTG));
PULLUP pullup1352 (.y(\~WR ));
PULLUP pullup1355 (.y(\op-T0-cmp ));
PULLUP pullup1356 (.y(net1356));
PULLUP pullup1357 (.y(net1357));
PULLUP pullup1358 (.y(net1358));
PULLUP pullup1364 (.y(net1364));
PULLUP pullup1368 (.y(net1368));
PULLUP pullup1369 (.y(net1369));
PULLUP pullup1370 (.y(Pout7));
PULLUP pullup1371 (.y(net1371));
PULLUP pullup1372 (.y(DC34));
PULLUP pullup1374 (.y(NMIL));
PULLUP pullup1375 (.y(net1375));
PULLUP pullup1376 (.y(net1376));
PULLUP pullup1377 (.y(net1377));
PULLUP pullup1379 (.y(net1379));
PULLUP pullup1380 (.y(net1380));
PULLUP pullup1381 (.y(\op-T3-jmp ));
PULLUP pullup1382 (.y(\brk-done ));
PULLUP pullup1383 (.y(net1383));
PULLUP pullup1384 (.y(ir2));
PULLUP pullup1385 (.y(\op-T5-mem-ind-idx ));
PULLUP pullup1386 (.y(net1386));
PULLUP pullup1389 (.y(net1389));
PULLUP pullup1391 (.y(net1391));
PULLUP pullup1392 (.y(net1392));
PULLUP pullup1394 (.y(notir5));
PULLUP pullup1396 (.y(\op-T0-shift-a ));
PULLUP pullup1398 (.y(\~(A+B)7 ));
PULLUP pullup1399 (.y(net1399));
PULLUP pullup1400 (.y(net1400));
PULLUP pullup1401 (.y(net1401));
PULLUP pullup1402 (.y(net1402));
PULLUP pullup1408 (.y(net1408));
PULLUP pullup1410 (.y(\pd7.clearIR ));
PULLUP pullup1412 (.y(net1412));
PULLUP pullup1413 (.y(net1413));
PULLUP pullup1414 (.y(alu3));
PULLUP pullup1415 (.y(dor6));
PULLUP pullup1416 (.y(net1416));
PULLUP pullup1419 (.y(\op-T0-cld/sed ));
PULLUP pullup1420 (.y(\op-T0-lda ));
PULLUP pullup1421 (.y(Pout2));
PULLUP pullup1423 (.y(net1423));
PULLUP pullup1425 (.y(\~C34 ));
PULLUP pullup1427 (.y(net1427));
PULLUP pullup1428 (.y(\op-T3-ind-x ));
PULLUP pullup1429 (.y(abh0));
PULLUP pullup1430 (.y(\x-op-T3-plp/pla ));
PULLUP pullup1433 (.y(net1433));
PULLUP pullup1434 (.y(notx1));
PULLUP pullup1439 (.y(noty6));
PULLUP pullup1440 (.y(net1440));
PULLUP pullup1441 (.y(net1441));
PULLUP pullup1444 (.y(Pout1));
PULLUP pullup1446 (.y(net1446));
PULLUP pullup1448 (.y(net1448));
PULLUP pullup1449 (.y(net1449));
PULLUP pullup1453 (.y(dor5));
PULLUP pullup1455 (.y(net1455));
PULLUP pullup1457 (.y(net1457));
PULLUP pullup1458 (.y(pclp6));
PULLUP pullup1459 (.y(\~(AxB)6 ));
PULLUP pullup1460 (.y(\pd6.clearIR ));
PULLUP pullup1462 (.y(net1462));
PULLUP pullup1463 (.y(net1463));
PULLUP pullup1464 (.y(net1464));
PULLUP pullup1465 (.y(VEC0));
PULLUP pullup1466 (.y(\op-rol/ror ));
PULLUP pullup1469 (.y(\~(AxB)5 ));
PULLUP pullup1471 (.y(net1471));
PULLUP pullup1474 (.y(net1474));
PULLUP pullup1475 (.y(dasb3));
PULLUP pullup1476 (.y(\x-op-T0-bit ));
PULLUP pullup1478 (.y(\op-T0-brk/rti ));
PULLUP pullup1481 (.y(VEC1));
PULLUP pullup1482 (.y(\op-T+-iny/dey ));
PULLUP pullup1484 (.y(noty2));
PULLUP pullup1486 (.y(net1486));
PULLUP pullup1487 (.y(\op-T3-plp/pla ));
PULLUP pullup1488 (.y(net1488));
PULLUP pullup1491 (.y(net1491));
PULLUP pullup1492 (.y(net1492));
PULLUP pullup1494 (.y(dasb7));
PULLUP pullup1495 (.y(net1495));
PULLUP pullup1496 (.y(pchp2));
PULLUP pullup1497 (.y(net1497));
PULLUP pullup1499 (.y(net1499));
PULLUP pullup1500 (.y(net1500));
PULLUP pullup1502 (.y(abl2));
PULLUP pullup1504 (.y(\op-T0-and ));
PULLUP pullup1506 (.y(\~C01 ));
PULLUP pullup1507 (.y(net1507));
PULLUP pullup1511 (.y(net1511));
PULLUP pullup1512 (.y(\op-T2-abs-y ));
PULLUP pullup1517 (.y(net1517));
PULLUP pullup1518 (.y(net1518));
PULLUP pullup1519 (.y(net1519));
PULLUP pullup1520 (.y(\op-plp/pla ));
PULLUP pullup1521 (.y(notx3));
PULLUP pullup1523 (.y(net1523));
PULLUP pullup1524 (.y(\op-T2-ind ));
PULLUP pullup1525 (.y(\~(AxB)0 ));
PULLUP pullup1526 (.y(net1526));
PULLUP pullup1531 (.y(net1531));
PULLUP pullup1534 (.y(net1534));
PULLUP pullup1540 (.y(\op-from-x ));
PULLUP pullup1541 (.y(net1541));
PULLUP pullup1542 (.y(net1542));
PULLUP pullup1543 (.y(\x-op-T0-txa ));
PULLUP pullup1544 (.y(BRtaken));
PULLUP pullup1548 (.y(net1548));
PULLUP pullup1549 (.y(net1549));
PULLUP pullup1552 (.y(net1552));
PULLUP pullup1557 (.y(\op-brk/rti ));
PULLUP pullup1560 (.y(net1560));
PULLUP pullup1561 (.y(notx7));
PULLUP pullup1562 (.y(\op-xy ));
PULLUP pullup1566 (.y(net1566));
PULLUP pullup1567 (.y(t3));
PULLUP pullup1569 (.y(\x-op-T4-rti ));
PULLUP pullup1571 (.y(\~C45 ));
PULLUP pullup1573 (.y(net1573));
PULLUP pullup1575 (.y(net1575));
PULLUP pullup1576 (.y(ir3));
PULLUP pullup1578 (.y(net1578));
PULLUP pullup1580 (.y(net1580));
PULLUP pullup1582 (.y(\op-T2-stack ));
PULLUP pullup1585 (.y(net1585));
PULLUP pullup1586 (.y(net1586));
PULLUP pullup1587 (.y(\pd3.clearIR ));
PULLUP pullup1588 (.y(net1588));
PULLUP pullup1589 (.y(\op-T4-jmp ));
PULLUP pullup1592 (.y(net1592));
PULLUP pullup1593 (.y(net1593));
PULLUP pullup1594 (.y(net1594));
PULLUP pullup1595 (.y(net1595));
PULLUP pullup1596 (.y(net1596));
PULLUP pullup1597 (.y(idl0));
PULLUP pullup1599 (.y(net1599));
PULLUP pullup1600 (.y(net1600));
PULLUP pullup1601 (.y(\op-sty/cpy-mem ));
PULLUP pullup1605 (.y(net1605));
PULLUP pullup1610 (.y(net1610));
PULLUP pullup1612 (.y(\op-T4-rts ));
PULLUP pullup1613 (.y(net1613));
PULLUP pullup1614 (.y(net1614));
PULLUP pullup1618 (.y(net1618));
PULLUP pullup1619 (.y(net1619));
PULLUP pullup1621 (.y(net1621));
PULLUP pullup1622 (.y(\pd0.clearIR ));
PULLUP pullup1623 (.y(\op-T0-eor ));
PULLUP pullup1626 (.y(ir1));
PULLUP pullup1628 (.y(\~A.B0 ));
PULLUP pullup1629 (.y(net1629));
PULLUP pullup1631 (.y(net1631));
PULLUP pullup1632 (.y(\~(A+B)5 ));
PULLUP pullup1634 (.y(dor2));
PULLUP pullup1635 (.y(net1635));
PULLUP pullup1637 (.y(alu2));
PULLUP pullup1638 (.y(net1638));
PULLUP pullup1640 (.y(noty7));
PULLUP pullup1641 (.y(net1641));
PULLUP pullup1642 (.y(net1642));
PULLUP pullup1643 (.y(net1643));
PULLUP pullup1646 (.y(\op-T+-bit ));
PULLUP pullup1647 (.y(pclp7));
PULLUP pullup1649 (.y(net1649));
PULLUP pullup1650 (.y(net1650));
PULLUP pullup1654 (.y(net1654));
PULLUP pullup1655 (.y(net1655));
PULLUP pullup1657 (.y(net1657));
PULLUP pullup1658 (.y(\op-T0-cpx/inx ));
PULLUP pullup1660 (.y(net1660));
PULLUP pullup1662 (.y(net1662));
PULLUP pullup1664 (.y(\op-T+-inx ));
PULLUP pullup1665 (.y(\op-T+-asl/rol-a ));
PULLUP pullup1668 (.y(net1668));
PULLUP pullup1671 (.y(\pd2.clearIR ));
PULLUP pullup1672 (.y(so));
PULLUP pullup1676 (.y(net1676));
PULLUP pullup1677 (.y(net1677));
PULLUP pullup1682 (.y(net1682));
PULLUP pullup1684 (.y(net1684));
PULLUP pullup1687 (.y(net1687));
PULLUP pullup1688 (.y(net1688));
PULLUP pullup1689 (.y(\op-EORS ));
PULLUP pullup1691 (.y(\~(A+B)2 ));
PULLUP pullup1694 (.y(net1694));
PULLUP pullup1697 (.y(net1697));
PULLUP pullup1704 (.y(dpc34_PCLC));
PULLUP pullup1705 (.y(net1705));
PULLUP pullup1708 (.y(\~op-T3-branch ));
PULLUP pullup1709 (.y(net1709));
PULLUP pullup1710 (.y(\op-T+-cpx/cpy-imm/zp ));
PULLUP pullup1711 (.y(net1711));
PULLUP pullup1712 (.y(net1712));
PULLUP pullup1714 (.y(net1714));
PULLUP pullup1715 (.y(net1715));
PULLUP pullup1716 (.y(net1716));
PULLUP pullup1717 (.y(net1717));
PULLUP pullup1718 (.y(net1718));
PULLUP pullup1719 (.y(net1719));
PULLUP pullup1720 (.y(net1720));
PULLUP pullup1721 (.y(\op-branch-done ));
PULLUP pullup1722 (.y(pchp0));
PULLUP pullup1724 (.y(net1724));

SW0 switch0 (.gate(pipeVectorA0), .cc(\0/ADL0 ));
SW1 switch1 (.gate(net1608), .cc(ab13));
SW0 switch2 (.gate(notalucout), .cc(alucout));
SW1 switch4 (.gate(net826), .cc(ab8));
SW0 switch5 (.gate(db1), .cc(net1319));
SW switch6 (.gate(\ADH/ABH ), .cc1(\~ABH6 ), .cc2(net1514));
SW0 switch8 (.gate(db2), .cc(net1199));
SW switch9 (.gate(cp1), .cc1(net524), .cc2(net1548));
SW0 switch10 (.gate(net190), .cc(net220));
SW1 switch11 (.gate(net38), .cc(net1247));
SW0 switch12 (.gate(alua1), .cc(net189));
SW0 switch13 (.gate(alua1), .cc(\~(A+B)1 ));
SW0 switch14 (.gate(cclk), .cc(net346));
SW1 switch15 (.gate(net1140), .cc(ab9));
SW0 switch16 (.gate(\op-from-x ), .cc(net508));
SW switch17 (.gate(cp1), .cc1(p0), .cc2(net1082));
SW switch18 (.gate(cp1), .cc1(net1451), .cc2(net212));
SW0 switch19 (.gate(net1247), .cc(dpc23_SBAC));
SW switch20 (.gate(cclk), .cc1(net1162), .cc2(net272));
SW switch21 (.gate(cclk), .cc1(net983), .cc2(nots0));
SW switch22 (.gate(notRdy0), .cc1(net1615), .cc2(net468));
SW switch23 (.gate(notRdy0), .cc1(net472), .cc2(net395));
SW switch24 (.gate(cp1), .cc1(net1495), .cc2(p3));
SW0 switch25 (.gate(abl0), .cc(net1100));
SW0 switch26 (.gate(abl0), .cc(net1660));
SW1 switch27 (.gate(abl0), .cc(net855));
SW0 switch28 (.gate(idb5), .cc(DBZ));
SW0 switch29 (.gate(pipeUNK05), .cc(net1616));
SW switch30 (.gate(C34), .cc1(\~(AxBxC)4 ), .cc2(net375));
SW0 switch31 (.gate(C34), .cc(\(AxB)4.~C34 ));
SW switch32 (.gate(cp1), .cc1(net928), .cc2(net1378));
SW switch33 (.gate(cp1), .cc1(net1309), .cc2(net74));
SW switch34 (.gate(cclk), .cc1(net518), .cc2(y6));
SW0 switch35 (.gate(p0), .cc(net31));
SW1 switch36 (.gate(cclk), .cc(dasb4));
SW switch37 (.gate(cclk), .cc1(net973), .cc2(nots4));
SW0 switch38 (.gate(net347), .cc(net510));
SW switch39 (.gate(cp1), .cc1(net1667), .cc2(net883));
SW0 switch40 (.gate(pipeT3out), .cc(net1456));
SW0 switch41 (.gate(\~op-branch-bit7 ), .cc(net307));
SW0 switch42 (.gate(\pd0.clearIR ), .cc(net409));
SW0 switch43 (.gate(net192), .cc(net25));
SW0 switch44 (.gate(notalu4), .cc(alu4));
SW switch45 (.gate(cclk), .cc1(y1), .cc2(net767));
SW switch46 (.gate(dpc11_SBADD), .cc1(sb1), .cc2(alua1));
SW switch47 (.gate(dpc11_SBADD), .cc1(sb2), .cc2(alua2));
SW switch48 (.gate(dpc11_SBADD), .cc1(alua3), .cc2(sb3));
SW switch49 (.gate(dpc11_SBADD), .cc1(alua4), .cc2(dasb4));
SW0 switch50 (.gate(RnWstretched), .cc(net794));
SW0 switch51 (.gate(RnWstretched), .cc(net794));
SW0 switch52 (.gate(net593), .cc(dpc4_SSB));
SW switch53 (.gate(dpc11_SBADD), .cc1(alua0), .cc2(dasb0));
SW switch54 (.gate(net600), .cc1(net613), .cc2(net1362));
SW switch55 (.gate(dpc11_SBADD), .cc1(alua5), .cc2(sb5));
SW switch56 (.gate(dpc11_SBADD), .cc1(alua6), .cc2(sb6));
SW0 switch57 (.gate(pch4), .cc(net1400));
SW switch58 (.gate(\~NMIG ), .cc1(net1092), .cc2(net480));
SW0 switch59 (.gate(\op-T2-stack ), .cc(net632));
SW0 switch60 (.gate(pch3), .cc(net923));
SW switch61 (.gate(\~C23 ), .cc1(\~(AxBxC)3 ), .cc2(net136));
SW0 switch62 (.gate(\~C23 ), .cc(\~(AxB3).C23 ));
SW switch63 (.gate(cclk), .cc1(net1347), .cc2(net1527));
SW0 switch64 (.gate(notalu6), .cc(alu6));
SW switch66 (.gate(net1457), .cc1(net1644), .cc2(net1495));
SW0 switch67 (.gate(notidl2), .cc(idl2));
SW0 switch68 (.gate(notidl2), .cc(idl2));
SW0 switch69 (.gate(notidl2), .cc(idl2));
SW0 switch70 (.gate(clearIR), .cc(\pd0.clearIR ));
SW0 switch71 (.gate(clearIR), .cc(\pd5.clearIR ));
SW switch72 (.gate(dpc1_SBY), .cc1(y6), .cc2(sb6));
SW switch73 (.gate(cp1), .cc1(net920), .cc2(net785));
SW0 switch74 (.gate(\~A.B7 ), .cc(net748));
SW1 switch75 (.gate(dpc14_SRS), .cc(\~aluresult7 ));
SW1 switch76 (.gate(net127), .cc(clk2out));
SW switch77 (.gate(dpc1_SBY), .cc1(y4), .cc2(dasb4));
SW0 switch78 (.gate(\op-lsr/ror/dec/inc ), .cc(net790));
SW0 switch79 (.gate(net763), .cc(dpc8_nDBADD));
SW0 switch80 (.gate(dor4), .cc(net147));
SW0 switch81 (.gate(dor4), .cc(net1463));
SW switch82 (.gate(H1x1), .cc1(Pout7), .cc2(idb7));
SW switch83 (.gate(H1x1), .cc1(idb2), .cc2(Pout2));
SW switch84 (.gate(cclk), .cc1(net513), .cc2(pipeUNK06));
SW switch85 (.gate(cclk), .cc1(net1673), .cc2(\op-T+-bit ));
SW switch86 (.gate(cclk), .cc1(net490), .cc2(notidl4));
SW0 switch87 (.gate(net311), .cc(net856));
SW0 switch88 (.gate(net311), .cc(net835));
SW0 switch89 (.gate(net783), .cc(net1158));
SW0 switch90 (.gate(net783), .cc(dpc34_PCLC));
SW0 switch91 (.gate(net783), .cc(net1253));
SW0 switch92 (.gate(net381), .cc(ab8));
SW0 switch93 (.gate(net381), .cc(ab8));
SW0 switch94 (.gate(net381), .cc(ab8));
SW0 switch95 (.gate(net381), .cc(ab8));
SW0 switch96 (.gate(net381), .cc(ab8));
SW0 switch97 (.gate(net381), .cc(ab8));
SW0 switch98 (.gate(net381), .cc(ab8));
SW0 switch99 (.gate(net152), .cc(net1343));
SW0 switch100 (.gate(\(AxB)0.~C0in ), .cc(\~(AxBxC)0 ));
SW0 switch101 (.gate(net810), .cc(net207));
SW0 switch102 (.gate(net819), .cc(net501));
SW0 switch103 (.gate(y1), .cc(noty1));
SW1 switch104 (.gate(net963), .cc(ab14));
SW0 switch105 (.gate(nnT2BR), .cc(net202));
SW0 switch106 (.gate(\~(A+B)2 ), .cc(net972));
SW0 switch107 (.gate(\op-T0-acc ), .cc(net1563));
SW0 switch108 (.gate(\op-T+-dex ), .cc(net844));
SW1 switch109 (.gate(abh3), .cc(net1296));
SW0 switch110 (.gate(abh3), .cc(net1346));
SW0 switch111 (.gate(abh3), .cc(net359));
SW0 switch112 (.gate(dpc12_0ADD), .cc(alua3));
SW0 switch113 (.gate(\pd7.clearIR ), .cc(\PD-0xx0xx0x ));
SW0 switch114 (.gate(\op-T0-ora ), .cc(net1145));
SW0 switch115 (.gate(notdor1), .cc(dor1));
SW switch116 (.gate(net1610), .cc1(net972), .cc2(DC34));
SW switch117 (.gate(cp1), .cc1(net653), .cc2(net1497));
SW0 switch118 (.gate(\~ABH7 ), .cc(abh7));
SW0 switch119 (.gate(net467), .cc(net10));
SW0 switch120 (.gate(net460), .cc(net692));
SW0 switch121 (.gate(\~pclp7 ), .cc(pclp7));
SW0 switch122 (.gate(net917), .cc(net1358));
SW switch123 (.gate(\ADH/ABH ), .cc1(\~ABH7 ), .cc2(net514));
SW0 switch124 (.gate(DBZ), .cc(\~DBZ ));
SW switch125 (.gate(cp1), .cc1(\short-circuit-branch-add ), .cc2(net1570));
SW switch126 (.gate(cclk), .cc1(net1179), .cc2(net393));
SW switch127 (.gate(dpc4_SSB), .cc1(net998), .cc2(sb3));
SW switch128 (.gate(dpc4_SSB), .cc1(net1389), .cc2(sb2));
SW0 switch129 (.gate(net1369), .cc(net1462));
SW1 switch130 (.gate(net1369), .cc(dpc38_PCLADL));
SW0 switch131 (.gate(\~op-store ), .cc(net816));
SW switch132 (.gate(dpc4_SSB), .cc1(net721), .cc2(sb7));
SW switch133 (.gate(dpc4_SSB), .cc1(net618), .cc2(sb6));
SW0 switch134 (.gate(net818), .cc(net1043));
SW1 switch135 (.gate(net818), .cc(dpc40_ADLPCL));
SW switch136 (.gate(dpc4_SSB), .cc1(net3), .cc2(dasb4));
SW0 switch137 (.gate(net270), .cc(net1426));
SW switch138 (.gate(alub5), .cc1(\~A.B5 ), .cc2(net1559));
SW0 switch139 (.gate(alub5), .cc(\~(A+B)5 ));
SW switch140 (.gate(cp1), .cc1(net1590), .cc2(net1083));
SW0 switch141 (.gate(x5), .cc(notx5));
SW switch142 (.gate(cp1), .cc1(net1424), .cc2(idl2));
SW0 switch143 (.gate(\op-T0-lda ), .cc(net1455));
SW0 switch144 (.gate(\op-T0-lda ), .cc(net397));
SW0 switch145 (.gate(idb7), .cc(net789));
SW0 switch146 (.gate(AxB3), .cc(\~(AxB)3 ));
SW0 switch147 (.gate(idb0), .cc(net624));
SW0 switch148 (.gate(net154), .cc(net75));
SW1 switch149 (.gate(net154), .cc(dpc20_ADDSB06));
SW0 switch150 (.gate(\op-T0-sbc ), .cc(net605));
SW0 switch151 (.gate(net1247), .cc(dpc1_SBY));
SW0 switch152 (.gate(\op-T2-stack ), .cc(net604));
SW0 switch153 (.gate(pch0), .cc(net1010));
SW1 switch154 (.gate(net798), .cc(db1));
SW1 switch155 (.gate(net798), .cc(db1));
SW0 switch156 (.gate(net453), .cc(net1264));
SW0 switch157 (.gate(\~ABL7 ), .cc(abl7));
SW0 switch158 (.gate(adl6), .cc(net1548));
SW0 switch159 (.gate(\op-T2-zp/zp-idx ), .cc(net1225));
SW0 switch160 (.gate(\~VEC ), .cc(net70));
SW0 switch161 (.gate(pipeT3out), .cc(net1366));
SW0 switch162 (.gate(net272), .cc(net952));
SW0 switch163 (.gate(net715), .cc(net426));
SW0 switch164 (.gate(net715), .cc(net914));
SW switch165 (.gate(net761), .cc1(net711), .cc2(net739));
SW1 switch166 (.gate(net1296), .cc(ab11));
SW1 switch167 (.gate(dor5), .cc(net373));
SW0 switch168 (.gate(net1312), .cc(\~NMIG ));
SW0 switch169 (.gate(net646), .cc(net812));
SW switch170 (.gate(cclk), .cc1(\~ABL5 ), .cc2(net210));
SW switch171 (.gate(\dpc36_~IPC ), .cc1(net1500), .cc2(net1706));
SW0 switch172 (.gate(\dpc36_~IPC ), .cc(net1345));
SW switch173 (.gate(net813), .cc1(net1101), .cc2(net1508));
SW0 switch174 (.gate(\op-T0-tay ), .cc(net11));
SW0 switch175 (.gate(net819), .cc(net1380));
SW1 switch176 (.gate(net714), .cc(dpc19_ADDSB7));
SW0 switch177 (.gate(net43), .cc(net818));
SW0 switch178 (.gate(\op-plp/pla ), .cc(net1107));
SW0 switch179 (.gate(net1002), .cc(net1130));
SW switch180 (.gate(cclk), .cc1(net779), .cc2(net805));
SW switch181 (.gate(cp1), .cc1(net1141), .cc2(net101));
SW switch182 (.gate(cclk), .cc1(net408), .cc2(notaluvout));
SW switch183 (.gate(net1581), .cc1(net1480), .cc2(\dpc36_~IPC ));
SW0 switch184 (.gate(net347), .cc(net191));
SW0 switch185 (.gate(notidl6), .cc(idl6));
SW0 switch186 (.gate(notidl6), .cc(idl6));
SW0 switch187 (.gate(notidl6), .cc(idl6));
SW0 switch188 (.gate(net1624), .cc(net169));
SW0 switch189 (.gate(net408), .cc(aluvout));
SW0 switch190 (.gate(ir3), .cc(notir3));
SW switch191 (.gate(cclk), .cc1(net1609), .cc2(notir5));
SW0 switch192 (.gate(pch7), .cc(net453));
SW0 switch193 (.gate(\op-T2-jmp-abs ), .cc(net368));
SW switch194 (.gate(BRtaken), .cc1(net405), .cc2(net1172));
SW0 switch195 (.gate(net1720), .cc(net373));
SW1 switch196 (.gate(net1720), .cc(net612));
SW1 switch197 (.gate(dor4), .cc(net1076));
SW0 switch198 (.gate(net646), .cc(net773));
SW0 switch199 (.gate(net982), .cc(net1141));
SW0 switch200 (.gate(net1135), .cc(net1203));
SW0 switch201 (.gate(net1135), .cc(net1629));
SW0 switch202 (.gate(net1258), .cc(net813));
SW0 switch203 (.gate(notRdy0), .cc(net720));
SW0 switch204 (.gate(net1045), .cc(net1371));
SW0 switch205 (.gate(net999), .cc(ab12));
SW0 switch206 (.gate(net999), .cc(ab12));
SW0 switch207 (.gate(net999), .cc(ab12));
SW0 switch208 (.gate(net999), .cc(ab12));
SW0 switch209 (.gate(net999), .cc(ab12));
SW0 switch210 (.gate(net999), .cc(ab12));
SW0 switch211 (.gate(net999), .cc(ab12));
SW switch212 (.gate(cclk), .cc1(pipeUNK22), .cc2(net29));
SW0 switch213 (.gate(net867), .cc(net876));
SW0 switch214 (.gate(\x-op-T0-tya ), .cc(net1717));
SW0 switch215 (.gate(alucout), .cc(\~alucout ));
SW0 switch216 (.gate(\op-T0-dex ), .cc(net1106));
SW0 switch217 (.gate(net241), .cc(net1033));
SW1 switch218 (.gate(net241), .cc(dpc21_ADDADL));
SW switch219 (.gate(net995), .cc1(net975), .cc2(net886));
SW0 switch220 (.gate(net201), .cc(net1371));
SW0 switch221 (.gate(\op-T2-abs-access ), .cc(net272));
SW0 switch222 (.gate(net846), .cc(net307));
SW switch223 (.gate(fetch), .cc1(net1183), .cc2(net541));
SW0 switch224 (.gate(D1x1), .cc(net380));
SW0 switch225 (.gate(net1061), .cc(\~pchp3 ));
SW switch226 (.gate(dpc7_SS), .cc1(net332), .cc2(s0));
SW1 switch227 (.gate(cclk), .cc(idb0));
SW0 switch228 (.gate(net621), .cc(net355));
SW0 switch229 (.gate(\~DBE ), .cc(net251));
SW0 switch230 (.gate(net1606), .cc(net188));
SW switch231 (.gate(\dpc42_DL/ADH ), .cc1(adh0), .cc2(net719));
SW switch232 (.gate(\dpc42_DL/ADH ), .cc1(adh1), .cc2(net87));
SW switch233 (.gate(\dpc42_DL/ADH ), .cc1(adh2), .cc2(net1424));
SW switch234 (.gate(\dpc42_DL/ADH ), .cc1(adh3), .cc2(net1661));
SW switch235 (.gate(\dpc42_DL/ADH ), .cc1(adh4), .cc2(net1095));
SW switch236 (.gate(\dpc42_DL/ADH ), .cc1(adh5), .cc2(net1387));
SW switch237 (.gate(\dpc42_DL/ADH ), .cc1(adh6), .cc2(net1014));
SW switch238 (.gate(\dpc42_DL/ADH ), .cc1(adh7), .cc2(net1147));
SW0 switch239 (.gate(\op-T5-brk ), .cc(net689));
SW0 switch240 (.gate(net805), .cc(net1534));
SW switch241 (.gate(cclk), .cc1(net326), .cc2(a6));
SW switch242 (.gate(cclk), .cc1(net1117), .cc2(pipeVectorA1));
SW switch243 (.gate(cp1), .cc1(net797), .cc2(notdor4));
SW0 switch244 (.gate(\brk-done ), .cc(net1087));
SW0 switch245 (.gate(pipeUNK32), .cc(net1178));
SW switch246 (.gate(alub0), .cc1(\~A.B0 ), .cc2(net316));
SW0 switch247 (.gate(alub0), .cc(\~(A+B)0 ));
SW switch248 (.gate(dpc6_SBS), .cc1(s5), .cc2(sb5));
SW switch249 (.gate(dpc6_SBS), .cc1(s6), .cc2(sb6));
SW switch250 (.gate(dpc6_SBS), .cc1(s3), .cc2(sb3));
SW switch251 (.gate(dpc6_SBS), .cc1(dasb4), .cc2(s4));
SW switch252 (.gate(dpc6_SBS), .cc1(s1), .cc2(sb1));
SW switch253 (.gate(dpc6_SBS), .cc1(s2), .cc2(sb2));
SW0 switch254 (.gate(net781), .cc(net802));
SW0 switch255 (.gate(\~(AxB)0 ), .cc(net406));
SW0 switch256 (.gate(\~(AxB)0 ), .cc(\(AxB)0.~C0in ));
SW0 switch257 (.gate(net647), .cc(\~C56 ));
SW0 switch258 (.gate(DC34), .cc(\~C34 ));
SW switch259 (.gate(cclk), .cc1(net242), .cc2(x3));
SW switch260 (.gate(cp1), .cc1(net931), .cc2(net1674));
SW switch261 (.gate(cp1), .cc1(net1526), .cc2(net1450));
SW0 switch262 (.gate(\op-T0 ), .cc(net638));
SW0 switch263 (.gate(net512), .cc(net154));
SW0 switch264 (.gate(net1247), .cc(dpc6_SBS));
SW0 switch265 (.gate(net1427), .cc(net1448));
SW0 switch266 (.gate(net223), .cc(net1357));
SW0 switch267 (.gate(net1219), .cc(net1002));
SW switch268 (.gate(H1x1), .cc1(idb0), .cc2(Pout0));
SW switch269 (.gate(cclk), .cc1(net604), .cc2(net1477));
SW switch270 (.gate(\~alucout ), .cc1(net367), .cc2(net1082));
SW0 switch271 (.gate(net265), .cc(net818));
SW0 switch272 (.gate(net1575), .cc(t2));
SW switch273 (.gate(net105), .cc1(\~(AxBxC)0 ), .cc2(net406));
SW0 switch274 (.gate(net105), .cc(\(AxB)0.~C0in ));
SW0 switch275 (.gate(net631), .cc(net1323));
SW1 switch276 (.gate(net631), .cc(dpc37_PCLDB));
SW0 switch277 (.gate(net544), .cc(net267));
SW0 switch278 (.gate(\op-T+-iny/dey ), .cc(net616));
SW1 switch279 (.gate(cclk), .cc(adl4));
SW0 switch280 (.gate(net101), .cc(net1364));
SW0 switch281 (.gate(\op-T0-ldx/tax/tsx ), .cc(net844));
SW0 switch282 (.gate(net1262), .cc(net1151));
SW switch283 (.gate(dpc7_SS), .cc1(net618), .cc2(s6));
SW switch284 (.gate(dpc7_SS), .cc1(net280), .cc2(s5));
SW switch285 (.gate(dpc7_SS), .cc1(net3), .cc2(s4));
SW switch286 (.gate(dpc7_SS), .cc1(net998), .cc2(s3));
SW switch287 (.gate(dpc7_SS), .cc1(net1389), .cc2(s2));
SW switch288 (.gate(dpc7_SS), .cc1(net694), .cc2(s1));
SW0 switch289 (.gate(adh3), .cc(net883));
SW0 switch290 (.gate(\~ABL6 ), .cc(abl6));
SW0 switch291 (.gate(\op-T4-mem-abs-idx ), .cc(net347));
SW0 switch292 (.gate(net781), .cc(net553));
SW0 switch293 (.gate(net1413), .cc(dpc32_PCHADH));
SW0 switch294 (.gate(\op-jmp ), .cc(net1649));
SW0 switch295 (.gate(s6), .cc(net1187));
SW switch296 (.gate(cp1), .cc1(net719), .cc2(idl0));
SW0 switch297 (.gate(\pd7.clearIR ), .cc(net1605));
SW0 switch298 (.gate(net279), .cc(net455));
SW1 switch299 (.gate(cclk), .cc(adh0));
SW0 switch300 (.gate(notx6), .cc(net1724));
SW0 switch301 (.gate(net612), .cc(db5));
SW0 switch302 (.gate(net612), .cc(db5));
SW0 switch303 (.gate(net612), .cc(db5));
SW0 switch304 (.gate(net612), .cc(db5));
SW0 switch305 (.gate(net612), .cc(db5));
SW0 switch306 (.gate(net612), .cc(db5));
SW0 switch307 (.gate(net612), .cc(db5));
SW0 switch308 (.gate(net445), .cc(net317));
SW0 switch309 (.gate(net445), .cc(net417));
SW0 switch310 (.gate(net445), .cc(net417));
SW0 switch311 (.gate(cp1), .cc(net127));
SW0 switch312 (.gate(net445), .cc(sync));
SW0 switch313 (.gate(net445), .cc(sync));
SW0 switch314 (.gate(net445), .cc(sync));
SW0 switch315 (.gate(net445), .cc(sync));
SW0 switch316 (.gate(net445), .cc(sync));
SW0 switch317 (.gate(\~ABH2 ), .cc(abh2));
SW0 switch318 (.gate(\brk-done ), .cc(net1215));
SW0 switch319 (.gate(AxB5), .cc(net547));
SW0 switch320 (.gate(AxB5), .cc(\~(AxB5).C45 ));
SW switch321 (.gate(dpc21_ADDADL), .cc1(alu2), .cc2(adl2));
SW switch322 (.gate(dpc21_ADDADL), .cc1(adl1), .cc2(alu1));
SW switch323 (.gate(dpc21_ADDADL), .cc1(adl0), .cc2(alu0));
SW0 switch324 (.gate(\op-T5-rti ), .cc(net1464));
SW0 switch325 (.gate(RESP), .cc(net501));
SW0 switch326 (.gate(net1699), .cc(net913));
SW0 switch327 (.gate(\x-op-T3-abs-idx ), .cc(net261));
SW0 switch328 (.gate(AxB1), .cc(net388));
SW switch329 (.gate(dpc0_YSB), .cc1(net564), .cc2(dasb0));
SW0 switch330 (.gate(net347), .cc(net335));
SW0 switch331 (.gate(net1602), .cc(net1596));
SW0 switch332 (.gate(net182), .cc(net442));
SW1 switch333 (.gate(dor1), .cc(net798));
SW switch334 (.gate(cclk), .cc1(net261), .cc2(pipeUNK36));
SW switch335 (.gate(cp1), .cc1(net959), .cc2(net323));
SW switch336 (.gate(cp1), .cc1(net1183), .cc2(net1605));
SW switch337 (.gate(net1595), .cc1(net1181), .cc2(net793));
SW0 switch338 (.gate(\~pclp0 ), .cc(pclp0));
SW0 switch339 (.gate(\op-T5-rts ), .cc(net182));
SW0 switch340 (.gate(net1452), .cc(net861));
SW0 switch341 (.gate(\op-T0-adc/sbc ), .cc(net1000));
SW0 switch342 (.gate(\~op-T3-branch ), .cc(net1055));
SW0 switch343 (.gate(net1305), .cc(dpc17_SUMS));
SW0 switch344 (.gate(net525), .cc(net800));
SW1 switch345 (.gate(net525), .cc(dpc26_ACDB));
SW0 switch346 (.gate(net1130), .cc(net80));
SW0 switch347 (.gate(\op-T3-jmp ), .cc(net980));
SW0 switch348 (.gate(ir0), .cc(net1133));
SW0 switch349 (.gate(ir0), .cc(notir0));
SW0 switch350 (.gate(net66), .cc(ab1));
SW0 switch351 (.gate(net66), .cc(ab1));
SW0 switch352 (.gate(net66), .cc(ab1));
SW0 switch353 (.gate(net66), .cc(ab1));
SW0 switch354 (.gate(cclk), .cc(dpc30_ADHPCH));
SW0 switch355 (.gate(cclk), .cc(dpc31_PCHPCH));
SW0 switch356 (.gate(net1341), .cc(net600));
SW0 switch357 (.gate(\op-T2-jsr ), .cc(net300));
SW0 switch358 (.gate(idb0), .cc(net1224));
SW switch359 (.gate(net335), .cc1(net1303), .cc2(net1397));
SW0 switch360 (.gate(net253), .cc(net279));
SW0 switch361 (.gate(net253), .cc(net1692));
SW1 switch362 (.gate(net1129), .cc(cclk));
SW0 switch363 (.gate(net1333), .cc(net906));
SW0 switch365 (.gate(net1081), .cc(net605));
SW0 switch366 (.gate(pipeUNK01), .cc(net1198));
SW1 switch367 (.gate(net424), .cc(notRdy0));
SW0 switch368 (.gate(pipeUNK31), .cc(net1178));
SW0 switch369 (.gate(net198), .cc(notRdy0));
SW0 switch370 (.gate(net198), .cc(net424));
SW switch371 (.gate(net335), .cc1(net1717), .cc2(net1604));
SW switch372 (.gate(dpc10_ADLADD), .cc1(adl0), .cc2(alub0));
SW0 switch373 (.gate(RESG), .cc(net1054));
SW switch374 (.gate(dpc4_SSB), .cc1(net694), .cc2(sb1));
SW0 switch375 (.gate(net869), .cc(ab13));
SW0 switch376 (.gate(net869), .cc(ab13));
SW0 switch377 (.gate(net869), .cc(ab13));
SW0 switch378 (.gate(net869), .cc(ab13));
SW0 switch379 (.gate(net869), .cc(ab13));
SW0 switch380 (.gate(net869), .cc(ab13));
SW0 switch381 (.gate(net869), .cc(ab13));
SW1 switch382 (.gate(net1076), .cc(db4));
SW1 switch383 (.gate(net1076), .cc(db4));
SW0 switch384 (.gate(pcl7), .cc(net641));
SW switch385 (.gate(dpc4_SSB), .cc1(net280), .cc2(sb5));
SW0 switch386 (.gate(\op-ror ), .cc(net544));
SW switch387 (.gate(\DA-C45 ), .cc1(net757), .cc2(net939));
SW switch388 (.gate(notRdy0), .cc1(net1456), .cc2(net428));
SW switch389 (.gate(notRdy0), .cc1(net12), .cc2(net1091));
SW0 switch390 (.gate(notRdy0), .cc(net16));
SW0 switch391 (.gate(db1), .cc(net213));
SW0 switch392 (.gate(pipeVectorA1), .cc(\0/ADL1 ));
SW0 switch393 (.gate(nots5), .cc(net280));
SW switch394 (.gate(cclk), .cc1(net1654), .cc2(a3));
SW switch395 (.gate(\ADH/ABH ), .cc1(net705), .cc2(\~ABH0 ));
SW0 switch396 (.gate(net521), .cc(net6));
SW1 switch397 (.gate(net317), .cc(net417));
SW0 switch398 (.gate(dpc29_0ADH17), .cc(adh1));
SW0 switch399 (.gate(RnWstretched), .cc(net1076));
SW0 switch400 (.gate(RnWstretched), .cc(net1076));
SW0 switch401 (.gate(RnWstretched), .cc(net1463));
SW switch402 (.gate(cp1), .cc1(p2), .cc2(net845));
SW0 switch403 (.gate(net1109), .cc(net1358));
SW0 switch404 (.gate(db3), .cc(net1281));
SW0 switch405 (.gate(\~C56 ), .cc(C56));
SW switch406 (.gate(\~C56 ), .cc1(net112), .cc2(C67));
SW switch407 (.gate(cclk), .cc1(net878), .cc2(net462));
SW0 switch408 (.gate(net330), .cc(net807));
SW0 switch409 (.gate(net1258), .cc(net1716));
SW switch410 (.gate(dpc30_ADHPCH), .cc1(pch3), .cc2(adh3));
SW switch411 (.gate(dpc30_ADHPCH), .cc1(pch2), .cc2(adh2));
SW switch412 (.gate(dpc30_ADHPCH), .cc1(pch5), .cc2(adh5));
SW switch413 (.gate(dpc30_ADHPCH), .cc1(pch4), .cc2(adh4));
SW switch414 (.gate(dpc30_ADHPCH), .cc1(pch7), .cc2(adh7));
SW switch415 (.gate(dpc30_ADHPCH), .cc1(pch6), .cc2(adh6));
SW1 switch416 (.gate(cclk), .cc(sb6));
SW switch417 (.gate(cclk), .cc1(net1187), .cc2(nots6));
SW0 switch418 (.gate(idb5), .cc(net1383));
SW switch419 (.gate(\ADH/ABH ), .cc1(net1667), .cc2(\~ABH3 ));
SW switch420 (.gate(cclk), .cc1(net1090), .cc2(net1683));
SW0 switch421 (.gate(net762), .cc(net1018));
SW0 switch422 (.gate(net135), .cc(clk2out));
SW0 switch423 (.gate(net135), .cc(clk2out));
SW0 switch424 (.gate(net135), .cc(clk2out));
SW0 switch425 (.gate(net135), .cc(clk2out));
SW1 switch426 (.gate(cclk), .cc(adh4));
SW1 switch427 (.gate(cclk), .cc(adl5));
SW switch428 (.gate(net440), .cc1(net366), .cc2(net1012));
SW0 switch429 (.gate(\~ABH4 ), .cc(abh4));
SW0 switch430 (.gate(net1162), .cc(net21));
SW switch431 (.gate(cclk), .cc1(net474), .cc2(net15));
SW switch432 (.gate(dpc2_XSB), .cc1(net1169), .cc2(dasb0));
SW0 switch433 (.gate(net962), .cc(\~DBE ));
SW0 switch434 (.gate(net1523), .cc(net963));
SW1 switch435 (.gate(net1523), .cc(net635));
SW0 switch436 (.gate(net1260), .cc(net1413));
SW1 switch437 (.gate(net1260), .cc(dpc32_PCHADH));
SW0 switch438 (.gate(net220), .cc(net130));
SW1 switch439 (.gate(net220), .cc(\ADL/ABL ));
SW0 switch440 (.gate(net400), .cc(net102));
SW1 switch441 (.gate(net400), .cc(net1696));
SW0 switch442 (.gate(net834), .cc(net1696));
SW0 switch443 (.gate(net834), .cc(net400));
SW0 switch444 (.gate(x7), .cc(notx7));
SW0 switch445 (.gate(net604), .cc(net656));
SW1 switch446 (.gate(net1545), .cc(ab10));
SW0 switch447 (.gate(\op-shift-right ), .cc(net1012));
SW0 switch448 (.gate(dpc35_PCHC), .cc(net949));
SW0 switch449 (.gate(dpc35_PCHC), .cc(net1406));
SW switch450 (.gate(dpc9_DBADD), .cc1(alub0), .cc2(idb0));
SW switch451 (.gate(cp1), .cc1(net402), .cc2(notRnWprepad));
SW0 switch452 (.gate(net358), .cc(net1129));
SW0 switch453 (.gate(net358), .cc(net1129));
SW switch454 (.gate(cclk), .cc1(net1717), .cc2(net1113));
SW switch455 (.gate(dpc2_XSB), .cc1(net871), .cc2(sb7));
SW1 switch456 (.gate(cclk), .cc(adh1));
SW switch457 (.gate(cclk), .cc1(net568), .cc2(notidl5));
SW0 switch458 (.gate(abl3), .cc(net138));
SW0 switch459 (.gate(abl3), .cc(net990));
SW1 switch460 (.gate(abl3), .cc(net1041));
SW0 switch461 (.gate(pipeUNK11), .cc(net1214));
SW0 switch462 (.gate(net1655), .cc(net182));
SW0 switch463 (.gate(a6), .cc(net1356));
SW0 switch464 (.gate(net378), .cc(t5));
SW0 switch465 (.gate(net35), .cc(net71));
SW1 switch466 (.gate(net35), .cc(dpc7_SS));
SW0 switch467 (.gate(\pipe~T0 ), .cc(net1180));
SW0 switch468 (.gate(\pipe~T0 ), .cc(net964));
SW0 switch469 (.gate(\op-T0-sbc ), .cc(net1304));
SW0 switch470 (.gate(nnT2BR), .cc(net1347));
SW0 switch471 (.gate(nnT2BR), .cc(net104));
SW switch472 (.gate(cp1), .cc1(net571), .cc2(net343));
SW switch473 (.gate(cclk), .cc1(net207), .cc2(net1061));
SW switch474 (.gate(net980), .cc1(net473), .cc2(net1004));
SW0 switch475 (.gate(rdy), .cc(net958));
SW1 switch476 (.gate(net963), .cc(ab14));
SW0 switch477 (.gate(net1240), .cc(\dpc43_DL/DB ));
SW switch478 (.gate(cclk), .cc1(\DC78.phi2 ), .cc2(DC78));
SW0 switch479 (.gate(\(AxB)6.~C56 ), .cc(\~(AxBxC)6 ));
SW0 switch480 (.gate(net781), .cc(net1170));
SW1 switch481 (.gate(net670), .cc(net1417));
SW0 switch482 (.gate(net994), .cc(ab10));
SW0 switch483 (.gate(net994), .cc(ab10));
SW0 switch484 (.gate(net994), .cc(ab10));
SW0 switch485 (.gate(net994), .cc(ab10));
SW0 switch486 (.gate(net994), .cc(ab10));
SW0 switch487 (.gate(net994), .cc(ab10));
SW0 switch488 (.gate(net994), .cc(ab10));
SW0 switch489 (.gate(noty6), .cc(net518));
SW switch490 (.gate(dpc7_SS), .cc1(s7), .cc2(net721));
SW0 switch491 (.gate(adh6), .cc(net880));
SW0 switch492 (.gate(net670), .cc(net747));
SW0 switch493 (.gate(net1472), .cc(net1480));
SW0 switch494 (.gate(\pd3.clearIR ), .cc(\PD-1xx000x0 ));
SW0 switch495 (.gate(\pd3.clearIR ), .cc(net1083));
SW switch496 (.gate(\~A.B0 ), .cc1(C01), .cc2(net942));
SW0 switch497 (.gate(net506), .cc(net877));
SW switch498 (.gate(net824), .cc1(net1278), .cc2(net1642));
SW switch499 (.gate(dpc13_ORS), .cc1(\~aluresult6 ), .cc2(\~(A+B)6 ));
SW0 switch500 (.gate(\op-T0-shift-a ), .cc(net1347));
SW0 switch501 (.gate(net1676), .cc(net634));
SW1 switch502 (.gate(net1676), .cc(net86));
SW switch503 (.gate(cclk), .cc1(notir0), .cc2(net310));
SW0 switch504 (.gate(net118), .cc(net1092));
SW0 switch505 (.gate(pipeUNK21), .cc(net572));
SW0 switch506 (.gate(sb6), .cc(net61));
SW0 switch507 (.gate(net1100), .cc(ab0));
SW0 switch508 (.gate(net1100), .cc(ab0));
SW0 switch509 (.gate(net1100), .cc(ab0));
SW0 switch510 (.gate(\op-T2-jsr ), .cc(net383));
SW0 switch511 (.gate(\op-T0-cpx/cpy/inx/iny ), .cc(net1560));
SW0 switch512 (.gate(nots4), .cc(net3));
SW switch513 (.gate(pipeUNK06), .cc1(net1422), .cc2(net754));
SW0 switch514 (.gate(pipeUNK06), .cc(net755));
SW switch515 (.gate(cclk), .cc1(net496), .cc2(nots5));
SW0 switch516 (.gate(net1223), .cc(net225));
SW1 switch517 (.gate(net1223), .cc(dpc9_DBADD));
SW0 switch518 (.gate(ir6), .cc(notir6));
SW0 switch519 (.gate(net1225), .cc(net1222));
SW switch520 (.gate(cp1), .cc1(net87), .cc2(idl1));
SW switch521 (.gate(dpc21_ADDADL), .cc1(adl3), .cc2(alu3));
SW switch522 (.gate(dpc21_ADDADL), .cc1(adl4), .cc2(alu4));
SW switch523 (.gate(cclk), .cc1(net844), .cc2(net459));
SW0 switch524 (.gate(db5), .cc(net568));
SW0 switch525 (.gate(net1517), .cc(net916));
SW switch526 (.gate(dpc21_ADDADL), .cc1(alu7), .cc2(adl7));
SW switch527 (.gate(dpc21_ADDADL), .cc1(adl5), .cc2(alu5));
SW switch528 (.gate(dpc21_ADDADL), .cc1(adl6), .cc2(alu6));
SW switch529 (.gate(net293), .cc1(net1402), .cc2(net57));
SW switch530 (.gate(net293), .cc1(net207), .cc2(net356));
SW0 switch531 (.gate(net293), .cc(net810));
SW switch532 (.gate(net335), .cc1(net734), .cc2(net1106));
SW0 switch533 (.gate(net807), .cc(net330));
SW0 switch534 (.gate(net990), .cc(net1041));
SW1 switch535 (.gate(net990), .cc(net138));
SW0 switch536 (.gate(net1357), .cc(net1575));
SW0 switch537 (.gate(net1097), .cc(dasb3));
SW switch538 (.gate(dpc13_ORS), .cc1(\~aluresult2 ), .cc2(\~(A+B)2 ));
SW switch539 (.gate(\op-T0-sbc ), .cc1(net51), .cc2(net29));
SW0 switch540 (.gate(net1635), .cc(dpc29_0ADH17));
SW switch541 (.gate(cp1), .cc1(net1641), .cc2(net237));
SW switch542 (.gate(cp1), .cc1(net724), .cc2(net409));
SW switch543 (.gate(net1662), .cc1(net1426), .cc2(net845));
SW0 switch544 (.gate(net267), .cc(net80));
SW switch545 (.gate(\~alucout ), .cc1(net387), .cc2(net916));
SW switch546 (.gate(dpc13_ORS), .cc1(\~(A+B)3 ), .cc2(\~aluresult3 ));
SW switch547 (.gate(C12), .cc1(\~(AxBxC)2 ), .cc2(net1572));
SW0 switch548 (.gate(C12), .cc(\(AxB)2.~C12 ));
SW switch549 (.gate(cclk), .cc1(\~aluresult3 ), .cc2(notalu3));
SW0 switch550 (.gate(net1109), .cc(net1130));
SW0 switch551 (.gate(net1417), .cc(clk1out));
SW0 switch552 (.gate(net1417), .cc(clk1out));
SW0 switch553 (.gate(net1417), .cc(clk1out));
SW0 switch554 (.gate(net1417), .cc(clk1out));
SW0 switch555 (.gate(net1417), .cc(clk1out));
SW switch556 (.gate(cclk), .cc1(net718), .cc2(notidl0));
SW0 switch557 (.gate(\A+B5 ), .cc(net165));
SW switch558 (.gate(net8), .cc1(net1584), .cc2(net345));
SW0 switch559 (.gate(dor2), .cc(net37));
SW0 switch560 (.gate(dor2), .cc(net224));
SW0 switch561 (.gate(net10), .cc(net176));
SW0 switch562 (.gate(net55), .cc(net628));
SW switch563 (.gate(net1614), .cc1(net299), .cc2(net1616));
SW0 switch564 (.gate(\~op-store ), .cc(net335));
SW0 switch565 (.gate(net664), .cc(net1697));
SW0 switch566 (.gate(VEC0), .cc(\~VEC ));
SW0 switch567 (.gate(\~(AxB)6 ), .cc(net122));
SW0 switch568 (.gate(\~(AxB)6 ), .cc(net1030));
SW0 switch569 (.gate(net772), .cc(net1305));
SW1 switch570 (.gate(net772), .cc(dpc17_SUMS));
SW0 switch571 (.gate(s5), .cc(net496));
SW0 switch572 (.gate(\~pclp2 ), .cc(pclp2));
SW0 switch573 (.gate(cclk), .cc(dpc23_SBAC));
SW0 switch574 (.gate(net459), .cc(net625));
SW0 switch575 (.gate(net43), .cc(net830));
SW switch577 (.gate(net755), .cc1(net566), .cc2(net580));
SW1 switch578 (.gate(dor2), .cc(net520));
SW0 switch579 (.gate(net732), .cc(net17));
SW0 switch580 (.gate(net732), .cc(clock1));
SW switch581 (.gate(cp1), .cc1(notRdy0), .cc2(net1679));
SW switch582 (.gate(cp1), .cc1(net223), .cc2(net1215));
SW0 switch583 (.gate(net748), .cc(\~C78 ));
SW0 switch584 (.gate(pipeUNK17), .cc(net511));
SW switch585 (.gate(\dpc43_DL/DB ), .cc1(idb0), .cc2(net719));
SW switch586 (.gate(\dpc43_DL/DB ), .cc1(idb1), .cc2(net87));
SW switch587 (.gate(\dpc43_DL/DB ), .cc1(idb2), .cc2(net1424));
SW switch588 (.gate(\dpc43_DL/DB ), .cc1(idb3), .cc2(net1661));
SW switch589 (.gate(\dpc43_DL/DB ), .cc1(idb4), .cc2(net1095));
SW switch590 (.gate(\dpc43_DL/DB ), .cc1(idb5), .cc2(net1387));
SW switch591 (.gate(\dpc43_DL/DB ), .cc1(idb6), .cc2(net1014));
SW switch592 (.gate(\dpc43_DL/DB ), .cc1(idb7), .cc2(net1147));
SW0 switch593 (.gate(NMIL), .cc(net1368));
SW1 switch594 (.gate(net322), .cc(ab7));
SW1 switch595 (.gate(net322), .cc(ab7));
SW1 switch596 (.gate(net322), .cc(ab7));
SW1 switch597 (.gate(net322), .cc(ab7));
SW0 switch598 (.gate(clock1), .cc(\op-T0-cpy/iny ));
SW0 switch599 (.gate(clock1), .cc(\op-T0-tay/ldy-not-idx ));
SW0 switch600 (.gate(clock1), .cc(\op-T0-iny/dey ));
SW0 switch601 (.gate(clock1), .cc(\x-op-T0-tya ));
SW0 switch602 (.gate(clock1), .cc(\x-op-T0-txa ));
SW0 switch603 (.gate(clock1), .cc(\op-T0-dex ));
SW0 switch604 (.gate(clock1), .cc(\op-T0-cpx/inx ));
SW0 switch605 (.gate(clock1), .cc(\op-T0-txs ));
SW0 switch606 (.gate(clock1), .cc(\op-T0-ldx/tax/tsx ));
SW0 switch607 (.gate(clock1), .cc(\op-T0-tsx ));
SW0 switch608 (.gate(clock1), .cc(\op-T0-ldy-mem ));
SW0 switch609 (.gate(clock1), .cc(\op-T0-jsr ));
SW0 switch610 (.gate(clock1), .cc(\op-T0-php/pha ));
SW0 switch611 (.gate(clock1), .cc(\op-T0-eor ));
SW0 switch612 (.gate(clock1), .cc(\op-T0-ora ));
SW0 switch613 (.gate(clock1), .cc(\op-T0 ));
SW0 switch614 (.gate(clock1), .cc(\op-T0-cpx/cpy/inx/iny ));
SW0 switch615 (.gate(clock1), .cc(\op-T0-cmp ));
SW0 switch616 (.gate(clock1), .cc(\op-T0-sbc ));
SW0 switch617 (.gate(clock1), .cc(\op-T0-adc/sbc ));
SW0 switch618 (.gate(clock1), .cc(\op-T0-tya ));
SW0 switch619 (.gate(clock1), .cc(\op-T0-txa ));
SW0 switch620 (.gate(clock1), .cc(\op-T0-pla ));
SW0 switch621 (.gate(clock1), .cc(\op-T0-lda ));
SW0 switch622 (.gate(clock1), .cc(\op-T0-acc ));
SW0 switch623 (.gate(clock1), .cc(\op-T0-tay ));
SW0 switch624 (.gate(clock1), .cc(\op-T0-shift-a ));
SW0 switch625 (.gate(clock1), .cc(\op-T0-tax ));
SW0 switch626 (.gate(clock1), .cc(\op-T0-bit ));
SW0 switch627 (.gate(clock1), .cc(\op-T0-and ));
SW0 switch628 (.gate(clock1), .cc(\op-branch-done ));
SW0 switch629 (.gate(clock1), .cc(\op-T0-shift-right-a ));
SW0 switch630 (.gate(clock1), .cc(\op-T0-brk/rti ));
SW0 switch631 (.gate(clock1), .cc(\op-T0-jmp ));
SW0 switch632 (.gate(clock1), .cc(\op-T0-cli/sei ));
SW0 switch633 (.gate(clock1), .cc(\op-T0-clc/sec ));
SW0 switch634 (.gate(clock1), .cc(\x-op-T0-bit ));
SW0 switch635 (.gate(clock1), .cc(\op-T0-plp ));
SW0 switch636 (.gate(clock1), .cc(\op-T0-cld/sed ));
SW switch637 (.gate(cclk), .cc1(y2), .cc2(net1491));
SW0 switch638 (.gate(net236), .cc(net272));
SW0 switch639 (.gate(net587), .cc(net299));
SW0 switch640 (.gate(ir6), .cc(\op-rol/ror ));
SW0 switch641 (.gate(ir6), .cc(\op-sty/cpy-mem ));
SW0 switch642 (.gate(ir6), .cc(\x-op-T0-tya ));
SW0 switch643 (.gate(ir6), .cc(\op-xy ));
SW0 switch644 (.gate(ir6), .cc(\x-op-T0-txa ));
SW0 switch645 (.gate(ir6), .cc(\op-from-x ));
SW0 switch646 (.gate(ir6), .cc(\op-T0-txs ));
SW0 switch647 (.gate(ir6), .cc(\op-T0-ldx/tax/tsx ));
SW0 switch648 (.gate(ir6), .cc(\op-T0-tsx ));
SW0 switch649 (.gate(ir6), .cc(\op-T0-ldy-mem ));
SW0 switch650 (.gate(ir6), .cc(\op-T0-tay/ldy-not-idx ));
SW0 switch651 (.gate(ir6), .cc(\op-T0-jsr ));
SW0 switch652 (.gate(ir6), .cc(\op-T5-brk ));
SW0 switch653 (.gate(ir6), .cc(\op-T0-ora ));
SW0 switch654 (.gate(ir6), .cc(\op-T4-brk/jsr ));
SW0 switch655 (.gate(ir6), .cc(\op-T2-jsr ));
SW0 switch656 (.gate(ir6), .cc(\op-shift ));
SW0 switch657 (.gate(ir6), .cc(\op-T5-jsr ));
SW0 switch658 (.gate(ir6), .cc(\op-T0-tya ));
SW0 switch659 (.gate(ir6), .cc(\op-T0-txa ));
SW0 switch660 (.gate(ir6), .cc(\op-T0-lda ));
SW0 switch661 (.gate(ir6), .cc(\op-T0-tay ));
SW0 switch662 (.gate(ir6), .cc(\op-T0-tax ));
SW0 switch663 (.gate(ir6), .cc(\op-T0-bit ));
SW0 switch664 (.gate(ir6), .cc(\op-T0-and ));
SW0 switch665 (.gate(ir6), .cc(\op-T2-brk ));
SW0 switch666 (.gate(ir6), .cc(\op-T3-jsr ));
SW0 switch667 (.gate(ir6), .cc(\op-sta/cmp ));
SW0 switch668 (.gate(ir6), .cc(\op-jsr ));
SW0 switch669 (.gate(ir6), .cc(\op-store ));
SW0 switch670 (.gate(ir6), .cc(\op-T4-brk ));
SW0 switch671 (.gate(ir6), .cc(\op-T2-php ));
SW0 switch672 (.gate(ir6), .cc(\xx-op-T5-jsr ));
SW0 switch673 (.gate(ir6), .cc(\op-asl/rol ));
SW0 switch674 (.gate(ir6), .cc(\op-T+-bit ));
SW0 switch675 (.gate(ir6), .cc(\op-T0-clc/sec ));
SW0 switch676 (.gate(ir6), .cc(\x-op-T0-bit ));
SW0 switch677 (.gate(ir6), .cc(\op-T0-plp ));
SW0 switch678 (.gate(ir6), .cc(\op-T+-asl/rol-a ));
SW0 switch679 (.gate(ir6), .cc(\~op-branch-bit6 ));
SW0 switch680 (.gate(ir6), .cc(\op-clv ));
SW switch681 (.gate(cclk), .cc1(net473), .cc2(pipeUNK33));
SW switch682 (.gate(cclk), .cc1(pipeUNK31), .cc2(net389));
SW0 switch683 (.gate(pcl3), .cc(net249));
SW switch684 (.gate(cclk), .cc1(pipeUNK32), .cc2(net1081));
SW0 switch685 (.gate(notRdy0), .cc(net1154));
SW0 switch686 (.gate(notRdy0), .cc(net180));
SW0 switch687 (.gate(net1202), .cc(net1367));
SW0 switch688 (.gate(net1202), .cc(net57));
SW0 switch689 (.gate(net307), .cc(net620));
SW0 switch690 (.gate(\op-T5-rti ), .cc(net256));
SW0 switch691 (.gate(pch6), .cc(net278));
SW0 switch692 (.gate(abl7), .cc(net171));
SW0 switch693 (.gate(abl7), .cc(net1026));
SW1 switch694 (.gate(abl7), .cc(net322));
SW0 switch695 (.gate(net551), .cc(net8));
SW switch696 (.gate(cclk), .cc1(net1620), .cc2(notir3));
SW0 switch698 (.gate(pipeUNK19), .cc(net1275));
SW0 switch699 (.gate(net491), .cc(dpc10_ADLADD));
SW0 switch700 (.gate(abl2), .cc(net642));
SW0 switch701 (.gate(abl2), .cc(net951));
SW1 switch702 (.gate(abl2), .cc(net1152));
SW0 switch703 (.gate(idb4), .cc(DBZ));
SW switch704 (.gate(net79), .cc1(net911), .cc2(net696));
SW switch705 (.gate(cclk), .cc1(\~aluresult5 ), .cc2(notalu5));
SW0 switch706 (.gate(notalucout), .cc(net1257));
SW switch707 (.gate(net1714), .cc1(net1189), .cc2(net262));
SW0 switch708 (.gate(AxB7), .cc(\~(AxB)7 ));
SW0 switch709 (.gate(idb6), .cc(net351));
SW0 switch710 (.gate(net43), .cc(net1541));
SW0 switch711 (.gate(net1529), .cc(net91));
SW0 switch712 (.gate(\op-T0-tax ), .cc(net11));
SW switch713 (.gate(cp1), .cc1(net854), .cc2(net1395));
SW0 switch714 (.gate(net1126), .cc(net1290));
SW switch715 (.gate(\~DA-ADD2 ), .cc1(net1556), .cc2(net986));
SW0 switch716 (.gate(\~DA-ADD2 ), .cc(net867));
SW0 switch717 (.gate(\op-T2-abs ), .cc(net1649));
SW0 switch718 (.gate(net1070), .cc(net1538));
SW0 switch719 (.gate(net1070), .cc(dpc35_PCHC));
SW0 switch720 (.gate(net1070), .cc(net200));
SW0 switch721 (.gate(ir4), .cc(\op-T0-iny/dey ));
SW0 switch722 (.gate(ir4), .cc(\op-T0-cpy/iny ));
SW0 switch723 (.gate(ir4), .cc(\op-T2-ind-x ));
SW0 switch724 (.gate(ir4), .cc(\x-op-T0-txa ));
SW0 switch725 (.gate(ir4), .cc(\op-T0-dex ));
SW0 switch726 (.gate(ir4), .cc(\op-T0-cpx/inx ));
SW0 switch727 (.gate(ir4), .cc(\op-T+-dex ));
SW0 switch728 (.gate(ir4), .cc(\op-T+-inx ));
SW0 switch729 (.gate(ir4), .cc(\op-T+-iny/dey ));
SW0 switch730 (.gate(ir4), .cc(\op-T0-tay/ldy-not-idx ));
SW0 switch731 (.gate(ir4), .cc(\op-T0-jsr ));
SW0 switch732 (.gate(ir4), .cc(\op-T5-brk ));
SW0 switch733 (.gate(ir4), .cc(\op-T0-php/pha ));
SW0 switch734 (.gate(ir4), .cc(\op-T4-rts ));
SW0 switch735 (.gate(ir4), .cc(\op-T3-plp/pla ));
SW0 switch736 (.gate(ir4), .cc(\op-T5-rti ));
SW0 switch737 (.gate(ir4), .cc(\op-jmp ));
SW0 switch738 (.gate(ir4), .cc(\op-T2-abs ));
SW0 switch739 (.gate(ir4), .cc(\op-T2-stack ));
SW0 switch740 (.gate(ir4), .cc(\op-T3-stack/bit/jmp ));
SW0 switch741 (.gate(ir4), .cc(\op-T4-brk/jsr ));
SW0 switch742 (.gate(ir4), .cc(\op-T4-rti ));
SW0 switch743 (.gate(ir4), .cc(\op-T3-ind-x ));
SW0 switch744 (.gate(ir4), .cc(\op-plp/pla ));
SW0 switch745 (.gate(ir4), .cc(\op-T4-ind-x ));
SW0 switch746 (.gate(ir4), .cc(\op-rti/rts ));
SW0 switch747 (.gate(ir4), .cc(\op-T2-jsr ));
SW0 switch748 (.gate(ir4), .cc(\op-T0-cpx/cpy/inx/iny ));
SW0 switch749 (.gate(ir4), .cc(\op-T3-jmp ));
SW0 switch750 (.gate(ir4), .cc(\op-T5-jsr ));
SW0 switch751 (.gate(ir4), .cc(\op-T2-stack-access ));
SW0 switch752 (.gate(ir4), .cc(\op-T+-shift-a ));
SW0 switch753 (.gate(ir4), .cc(\op-T0-txa ));
SW0 switch754 (.gate(ir4), .cc(\op-T0-pla ));
SW0 switch755 (.gate(ir4), .cc(\op-T0-tay ));
SW0 switch756 (.gate(ir4), .cc(\op-T0-shift-a ));
SW0 switch757 (.gate(ir4), .cc(\op-T0-tax ));
SW0 switch758 (.gate(ir4), .cc(\op-T0-bit ));
SW0 switch759 (.gate(ir4), .cc(\op-T2-pha ));
SW0 switch760 (.gate(ir4), .cc(\op-T0-shift-right-a ));
SW0 switch761 (.gate(ir4), .cc(\op-T2-brk ));
SW0 switch762 (.gate(ir4), .cc(\op-T3-jsr ));
SW0 switch763 (.gate(ir4), .cc(\op-T5-rts ));
SW0 switch764 (.gate(ir4), .cc(\op-T0-brk/rti ));
SW0 switch765 (.gate(ir4), .cc(\op-T0-jmp ));
SW0 switch766 (.gate(ir4), .cc(\op-T5-ind-x ));
SW0 switch767 (.gate(ir4), .cc(\op-brk/rti ));
SW0 switch768 (.gate(ir4), .cc(\op-jsr ));
SW0 switch769 (.gate(ir4), .cc(\x-op-jmp ));
SW0 switch770 (.gate(ir4), .cc(\op-push/pull ));
SW0 switch771 (.gate(ir4), .cc(\op-T4-brk ));
SW0 switch772 (.gate(ir4), .cc(\op-T2-php ));
SW0 switch773 (.gate(ir4), .cc(\op-T2-php/pha ));
SW0 switch774 (.gate(ir4), .cc(\op-T4-jmp ));
SW0 switch775 (.gate(ir4), .cc(\op-T5-rti/rts ));
SW0 switch776 (.gate(ir4), .cc(\xx-op-T5-jsr ));
SW0 switch777 (.gate(ir4), .cc(\op-T2-jmp-abs ));
SW0 switch778 (.gate(ir4), .cc(\x-op-T3-plp/pla ));
SW0 switch779 (.gate(ir4), .cc(\op-T+-bit ));
SW0 switch780 (.gate(ir4), .cc(\x-op-T0-bit ));
SW0 switch781 (.gate(ir4), .cc(\op-T0-plp ));
SW0 switch782 (.gate(ir4), .cc(\x-op-T4-rti ));
SW0 switch783 (.gate(ir4), .cc(\op-T+-cpx/cpy-abs ));
SW0 switch784 (.gate(ir4), .cc(\op-T+-asl/rol-a ));
SW0 switch785 (.gate(ir4), .cc(\op-T+-cpx/cpy-imm/zp ));
SW0 switch786 (.gate(ir4), .cc(\x-op-push/pull ));
SW0 switch787 (.gate(ir4), .cc(\op-T3-mem-abs ));
SW0 switch788 (.gate(ir4), .cc(\op-T2-mem-zp ));
SW0 switch789 (.gate(net1300), .cc(ir2));
SW switch790 (.gate(cp1), .cc1(net416), .cc2(net1016));
SW0 switch791 (.gate(notalu2), .cc(alu2));
SW switch792 (.gate(BRtaken), .cc1(net586), .cc2(net1330));
SW switch793 (.gate(BRtaken), .cc1(net586), .cc2(net1330));
SW switch794 (.gate(cclk), .cc1(pipeUNK14), .cc2(net318));
SW0 switch795 (.gate(ir7), .cc(\op-rol/ror ));
SW0 switch796 (.gate(ir7), .cc(\op-T0-jsr ));
SW0 switch797 (.gate(ir7), .cc(\op-T5-brk ));
SW0 switch798 (.gate(ir7), .cc(\op-T0-php/pha ));
SW0 switch799 (.gate(ir7), .cc(\op-T4-rts ));
SW0 switch800 (.gate(ir7), .cc(\op-T3-plp/pla ));
SW0 switch801 (.gate(ir7), .cc(\op-T5-rti ));
SW0 switch802 (.gate(ir7), .cc(\op-ror ));
SW0 switch803 (.gate(ir7), .cc(\op-T0-eor ));
SW0 switch804 (.gate(ir7), .cc(\op-jmp ));
SW0 switch805 (.gate(ir7), .cc(\op-T0-ora ));
SW0 switch806 (.gate(ir7), .cc(\op-T2-stack ));
SW0 switch807 (.gate(ir7), .cc(\op-T3-stack/bit/jmp ));
SW0 switch808 (.gate(ir7), .cc(\op-T4-brk/jsr ));
SW0 switch809 (.gate(ir7), .cc(\op-T4-rti ));
SW0 switch810 (.gate(ir7), .cc(\op-plp/pla ));
SW0 switch811 (.gate(ir7), .cc(\op-rti/rts ));
SW0 switch812 (.gate(ir7), .cc(\op-T2-jsr ));
SW0 switch813 (.gate(ir7), .cc(\op-T3-jmp ));
SW0 switch814 (.gate(ir7), .cc(\op-shift ));
SW0 switch815 (.gate(ir7), .cc(\op-T5-jsr ));
SW0 switch816 (.gate(ir7), .cc(\op-T2-stack-access ));
SW0 switch817 (.gate(ir7), .cc(\op-T+-ora/and/eor/adc ));
SW0 switch818 (.gate(ir7), .cc(\op-T+-shift-a ));
SW0 switch819 (.gate(ir7), .cc(\op-T0-pla ));
SW0 switch820 (.gate(ir7), .cc(\op-T0-shift-a ));
SW0 switch821 (.gate(ir7), .cc(\op-T0-bit ));
SW0 switch822 (.gate(ir7), .cc(\op-T0-and ));
SW0 switch823 (.gate(ir7), .cc(\op-T2-pha ));
SW0 switch824 (.gate(ir7), .cc(\op-T0-shift-right-a ));
SW0 switch825 (.gate(ir7), .cc(\op-shift-right ));
SW0 switch826 (.gate(ir7), .cc(\op-T2-brk ));
SW0 switch827 (.gate(ir7), .cc(\op-T3-jsr ));
SW0 switch828 (.gate(ir7), .cc(\op-T5-rts ));
SW0 switch829 (.gate(ir7), .cc(\op-T0-brk/rti ));
SW0 switch830 (.gate(ir7), .cc(\op-T0-jmp ));
SW0 switch831 (.gate(ir7), .cc(\op-brk/rti ));
SW0 switch832 (.gate(ir7), .cc(\op-jsr ));
SW0 switch833 (.gate(ir7), .cc(\x-op-jmp ));
SW0 switch834 (.gate(ir7), .cc(\op-push/pull ));
SW0 switch835 (.gate(ir7), .cc(\op-T4-brk ));
SW0 switch836 (.gate(ir7), .cc(\op-T2-php ));
SW0 switch837 (.gate(ir7), .cc(\op-T2-php/pha ));
SW0 switch838 (.gate(ir7), .cc(\op-T4-jmp ));
SW0 switch839 (.gate(ir7), .cc(\op-T5-rti/rts ));
SW0 switch840 (.gate(ir7), .cc(\xx-op-T5-jsr ));
SW0 switch841 (.gate(ir7), .cc(\op-T2-jmp-abs ));
SW0 switch842 (.gate(ir7), .cc(\x-op-T3-plp/pla ));
SW0 switch843 (.gate(ir7), .cc(\op-asl/rol ));
SW0 switch844 (.gate(ir7), .cc(\op-T0-cli/sei ));
SW0 switch845 (.gate(ir7), .cc(\op-T+-bit ));
SW0 switch846 (.gate(ir7), .cc(\op-T0-clc/sec ));
SW0 switch847 (.gate(ir7), .cc(\x-op-T0-bit ));
SW0 switch848 (.gate(ir7), .cc(\op-T0-plp ));
SW0 switch849 (.gate(ir7), .cc(\x-op-T4-rti ));
SW0 switch850 (.gate(ir7), .cc(\op-T+-asl/rol-a ));
SW0 switch851 (.gate(ir7), .cc(\x-op-push/pull ));
SW0 switch852 (.gate(ir7), .cc(\~op-branch-bit7 ));
SW0 switch853 (.gate(\~A.B4 ), .cc(net1310));
SW1 switch854 (.gate(net963), .cc(ab14));
SW0 switch855 (.gate(\~op-branch-bit6 ), .cc(net846));
SW0 switch856 (.gate(\pipe~WR.phi2 ), .cc(notRnWprepad));
SW switch857 (.gate(net243), .cc1(net566), .cc2(net802));
SW0 switch858 (.gate(\DA-AB2 ), .cc(\DA-AxB2 ));
SW0 switch859 (.gate(\DA-AB2 ), .cc(net1610));
SW0 switch860 (.gate(adl7), .cc(net1046));
SW0 switch861 (.gate(net1107), .cc(net389));
SW switch862 (.gate(\ADL/ABL ), .cc1(net416), .cc2(\~ABL1 ));
SW0 switch863 (.gate(net1007), .cc(dpc35_PCHC));
SW0 switch864 (.gate(net1673), .cc(net754));
SW switch865 (.gate(\ADL/ABL ), .cc1(net1636), .cc2(\~ABL2 ));
SW0 switch866 (.gate(y2), .cc(noty2));
SW0 switch867 (.gate(AxB7), .cc(net1013));
SW0 switch868 (.gate(AxB7), .cc(\~(AxB7).C67 ));
SW0 switch869 (.gate(net291), .cc(net1157));
SW1 switch870 (.gate(net291), .cc(\dpc41_DL/ADL ));
SW0 switch871 (.gate(\op-T2-ind ), .cc(net1225));
SW0 switch872 (.gate(\op-branch-done ), .cc(net10));
SW0 switch873 (.gate(net278), .cc(net1488));
SW0 switch874 (.gate(net462), .cc(net1278));
SW0 switch875 (.gate(net599), .cc(\dpc22_~DSA ));
SW0 switch876 (.gate(net692), .cc(net441));
SW1 switch877 (.gate(net692), .cc(dpc1_SBY));
SW0 switch878 (.gate(\op-T4-ind-x ), .cc(net300));
SW0 switch879 (.gate(net760), .cc(INTG));
SW0 switch880 (.gate(idb2), .cc(net458));
SW0 switch881 (.gate(\~pchp4 ), .cc(pchp4));
SW0 switch882 (.gate(net383), .cc(net917));
SW0 switch883 (.gate(pcl5), .cc(net386));
SW0 switch884 (.gate(notRdy0), .cc(net1649));
SW switch885 (.gate(net16), .cc1(net472), .cc2(net1366));
SW0 switch886 (.gate(pipeUNK18), .cc(net850));
SW0 switch887 (.gate(RnWstretched), .cc(net147));
SW0 switch888 (.gate(RnWstretched), .cc(net147));
SW0 switch889 (.gate(\op-T5-mem-ind-idx ), .cc(net347));
SW switch890 (.gate(cp1), .cc1(net1132), .cc2(net1087));
SW0 switch891 (.gate(notRdy0), .cc(net1180));
SW switch892 (.gate(cclk), .cc1(pipeT4out), .cc2(net188));
SW0 switch893 (.gate(\~(AxB5).C45 ), .cc(\~(AxBxC)5 ));
SW1 switch894 (.gate(abh6), .cc(net963));
SW0 switch895 (.gate(abh6), .cc(net1523));
SW0 switch896 (.gate(abh6), .cc(net635));
SW0 switch897 (.gate(net225), .cc(dpc9_DBADD));
SW0 switch898 (.gate(AxB3), .cc(net136));
SW0 switch899 (.gate(AxB3), .cc(\~(AxB3).C23 ));
SW0 switch900 (.gate(\~(A+B)1 ), .cc(\A+B1 ));
SW0 switch901 (.gate(\~(A+B)1 ), .cc(AxB1));
SW0 switch902 (.gate(net440), .cc(net1555));
SW0 switch903 (.gate(net432), .cc(net1686));
SW0 switch904 (.gate(net432), .cc(net1097));
SW0 switch905 (.gate(net635), .cc(ab14));
SW0 switch906 (.gate(net635), .cc(ab14));
SW0 switch907 (.gate(net635), .cc(ab14));
SW0 switch908 (.gate(net635), .cc(ab14));
SW0 switch909 (.gate(net635), .cc(ab14));
SW0 switch910 (.gate(net635), .cc(ab14));
SW0 switch911 (.gate(net635), .cc(ab14));
SW0 switch912 (.gate(net43), .cc(net1534));
SW0 switch913 (.gate(nnT2BR), .cc(net1330));
SW0 switch914 (.gate(nots7), .cc(net721));
SW switch915 (.gate(cclk), .cc1(net1225), .cc2(pipedpc28));
SW0 switch916 (.gate(net726), .cc(net630));
SW0 switch917 (.gate(net1195), .cc(net1191));
SW1 switch918 (.gate(net1195), .cc(net1254));
SW0 switch919 (.gate(\branch-back.phi1 ), .cc(net1055));
SW0 switch920 (.gate(net221), .cc(net251));
SW0 switch921 (.gate(net221), .cc(net251));
SW0 switch922 (.gate(notRdy0), .cc(net372));
SW switch923 (.gate(notRdy0), .cc1(net1365), .cc2(net1085));
SW switch924 (.gate(cclk), .cc1(net359), .cc2(\~ABH3 ));
SW switch925 (.gate(cp1), .cc1(\branch-back ), .cc2(net756));
SW switch926 (.gate(cp1), .cc1(net457), .cc2(notdor3));
SW0 switch927 (.gate(net255), .cc(dpc31_PCHPCH));
SW1 switch928 (.gate(net1140), .cc(ab9));
SW0 switch929 (.gate(notdor2), .cc(dor2));
SW0 switch930 (.gate(net383), .cc(net1040));
SW0 switch931 (.gate(net383), .cc(net1040));
SW0 switch932 (.gate(alu2), .cc(\~DA-ADD2 ));
SW switch933 (.gate(net270), .cc1(net1445), .cc2(net1495));
SW0 switch934 (.gate(net1593), .cc(net1552));
SW1 switch935 (.gate(net1593), .cc(dpc14_SRS));
SW switch936 (.gate(dpc16_EORS), .cc1(\~(AxB)0 ), .cc2(\~aluresult0 ));
SW switch937 (.gate(dpc16_EORS), .cc1(\~aluresult1 ), .cc2(\~(AxB)1 ));
SW switch938 (.gate(dpc16_EORS), .cc1(\~(AxB)2 ), .cc2(\~aluresult2 ));
SW switch939 (.gate(dpc16_EORS), .cc1(\~(AxB)3 ), .cc2(\~aluresult3 ));
SW switch940 (.gate(dpc16_EORS), .cc1(\~(AxB)4 ), .cc2(\~aluresult4 ));
SW switch941 (.gate(dpc16_EORS), .cc1(\~(AxB)5 ), .cc2(\~aluresult5 ));
SW switch942 (.gate(dpc16_EORS), .cc1(\~(AxB)6 ), .cc2(\~aluresult6 ));
SW switch943 (.gate(dpc16_EORS), .cc1(\~aluresult7 ), .cc2(\~(AxB)7 ));
SW0 switch944 (.gate(\op-T4 ), .cc(net256));
SW switch945 (.gate(net16), .cc1(net1558), .cc2(net428));
SW switch946 (.gate(\op-asl/rol ), .cc1(\~op-set-C ), .cc2(net591));
SW0 switch948 (.gate(Pout3), .cc(net1053));
SW0 switch949 (.gate(clock2), .cc(\op-T+-dex ));
SW0 switch950 (.gate(clock2), .cc(\op-T+-inx ));
SW0 switch951 (.gate(clock2), .cc(\op-T+-iny/dey ));
SW0 switch952 (.gate(clock2), .cc(\op-T+-ora/and/eor/adc ));
SW0 switch953 (.gate(clock2), .cc(\op-T+-adc/sbc ));
SW0 switch954 (.gate(clock2), .cc(\op-T+-shift-a ));
SW0 switch955 (.gate(clock2), .cc(\op-T+-bit ));
SW0 switch956 (.gate(clock2), .cc(\x-op-T+-adc/sbc ));
SW0 switch957 (.gate(clock2), .cc(\op-T+-cmp ));
SW0 switch958 (.gate(clock2), .cc(\op-T+-cpx/cpy-abs ));
SW0 switch959 (.gate(clock2), .cc(\op-T+-asl/rol-a ));
SW0 switch960 (.gate(clock2), .cc(\op-T+-cpx/cpy-imm/zp ));
SW1 switch961 (.gate(cclk), .cc(idb3));
SW switch962 (.gate(cclk), .cc1(net1694), .cc2(x2));
SW switch963 (.gate(dpc6_SBS), .cc1(dasb0), .cc2(s0));
SW0 switch964 (.gate(net1120), .cc(net137));
SW0 switch966 (.gate(idb6), .cc(DBZ));
SW0 switch967 (.gate(net368), .cc(net218));
SW switch968 (.gate(\DA-C01 ), .cc1(net319), .cc2(net1707));
SW0 switch969 (.gate(\DA-C01 ), .cc(net388));
SW0 switch970 (.gate(net1578), .cc(net1368));
SW0 switch971 (.gate(net1027), .cc(net476));
SW0 switch972 (.gate(\op-T4-jmp ), .cc(net368));
SW0 switch973 (.gate(\op-T4-jmp ), .cc(net104));
SW0 switch974 (.gate(\~ABL0 ), .cc(abl0));
SW0 switch975 (.gate(net440), .cc(\~WR ));
SW0 switch976 (.gate(net440), .cc(net104));
SW0 switch977 (.gate(net440), .cc(net812));
SW0 switch978 (.gate(net1585), .cc(net962));
SW0 switch979 (.gate(\~(A+B)7 ), .cc(net1489));
SW switch980 (.gate(\op-T2-idx-x-xy ), .cc1(net1103), .cc2(net1106));
SW0 switch981 (.gate(net979), .cc(net1347));
SW0 switch982 (.gate(\op-T5-brk ), .cc(net1464));
SW0 switch983 (.gate(pd2), .cc(\pd2.clearIR ));
SW0 switch984 (.gate(net1343), .cc(net911));
SW0 switch985 (.gate(net790), .cc(\op-rmw ));
SW0 switch986 (.gate(net1054), .cc(net70));
SW0 switch987 (.gate(\x-op-T0-txa ), .cc(net1106));
SW0 switch988 (.gate(sb1), .cc(net320));
SW switch989 (.gate(dpc37_PCLDB), .cc1(idb0), .cc2(pclp0));
SW1 switch990 (.gate(abh5), .cc(net1608));
SW0 switch991 (.gate(abh5), .cc(net1423));
SW0 switch992 (.gate(abh5), .cc(net869));
SW switch993 (.gate(dpc37_PCLDB), .cc1(idb2), .cc2(pclp2));
SW0 switch994 (.gate(\op-clv ), .cc(net340));
SW0 switch995 (.gate(notRdy0), .cc(\brk-done ));
SW switch996 (.gate(\op-T0-adc/sbc ), .cc1(net673), .cc2(net1053));
SW switch997 (.gate(fetch), .cc1(net703), .cc2(net927));
SW0 switch998 (.gate(net415), .cc(net931));
SW0 switch999 (.gate(net88), .cc(net1375));
SW0 switch1000 (.gate(\branch-forward.phi1 ), .cc(\branch-back.phi1 ));
SW switch1001 (.gate(\~C01 ), .cc1(\~(AxBxC)1 ), .cc2(net1388));
SW0 switch1002 (.gate(\~C01 ), .cc(\~(AxB1).C01 ));
SW0 switch1003 (.gate(RnWstretched), .cc(net7));
SW0 switch1004 (.gate(RnWstretched), .cc(net7));
SW0 switch1005 (.gate(RnWstretched), .cc(net466));
SW0 switch1006 (.gate(pipeUNK27), .cc(net920));
SW0 switch1007 (.gate(\(AxB)4.~C34 ), .cc(\~(AxBxC)4 ));
SW switch1008 (.gate(cp1), .cc1(notRdy0), .cc2(net902));
SW0 switch1009 (.gate(ir2), .cc(notir2));
SW switch1010 (.gate(cclk), .cc1(net1675), .cc2(notir6));
SW0 switch1011 (.gate(net25), .cc(net674));
SW switch1012 (.gate(cclk), .cc1(net1588), .cc2(pd5));
SW switch1013 (.gate(cclk), .cc1(pd3), .cc2(net1281));
SW switch1014 (.gate(cclk), .cc1(pd4), .cc2(net1075));
SW switch1015 (.gate(cclk), .cc1(net929), .cc2(a1));
SW0 switch1016 (.gate(net688), .cc(net1223));
SW switch1017 (.gate(cclk), .cc1(net1638), .cc2(notidl6));
SW switch1018 (.gate(\A+B2 ), .cc1(\~(AxB)2 ), .cc2(net716));
SW0 switch1019 (.gate(net510), .cc(net1716));
SW0 switch1020 (.gate(net1113), .cc(net161));
SW0 switch1021 (.gate(net861), .cc(\brk-done ));
SW0 switch1022 (.gate(net1247), .cc(dpc8_nDBADD));
SW switch1023 (.gate(net471), .cc1(db6), .cc2(db6));
SW0 switch1024 (.gate(net471), .cc(db6));
SW0 switch1025 (.gate(net471), .cc(db6));
SW0 switch1026 (.gate(net471), .cc(db6));
SW0 switch1027 (.gate(net471), .cc(db6));
SW0 switch1028 (.gate(net471), .cc(db6));
SW0 switch1029 (.gate(net471), .cc(db6));
SW0 switch1030 (.gate(net471), .cc(db6));
SW0 switch1031 (.gate(net471), .cc(db6));
SW0 switch1032 (.gate(RnWstretched), .cc(net1325));
SW0 switch1033 (.gate(RnWstretched), .cc(net1325));
SW0 switch1034 (.gate(RnWstretched), .cc(net769));
SW1 switch1035 (.gate(net358), .cc(net1467));
SW switch1036 (.gate(cp1), .cc1(net463), .cc2(net1094));
SW switch1037 (.gate(fetch), .cc1(net1590), .cc2(net1620));
SW0 switch1038 (.gate(net645), .cc(net1368));
SW0 switch1039 (.gate(notRdy0), .cc(net1275));
SW0 switch1040 (.gate(adh1), .cc(net1267));
SW switch1041 (.gate(cp1), .cc1(net494), .cc2(net514));
SW0 switch1042 (.gate(net954), .cc(net279));
SW0 switch1043 (.gate(net954), .cc(net367));
SW0 switch1044 (.gate(net236), .cc(net1427));
SW0 switch1045 (.gate(\op-T0-jsr ), .cc(net1464));
SW0 switch1046 (.gate(\~pchp2 ), .cc(pchp2));
SW switch1047 (.gate(cclk), .cc1(net1251), .cc2(y7));
SW0 switch1048 (.gate(adl4), .cc(net1519));
SW switch1049 (.gate(cp1), .cc1(net262), .cc2(net1447));
SW0 switch1050 (.gate(\op-ORS ), .cc(\op-SUMS ));
SW switch1051 (.gate(\ADL/ABL ), .cc1(net246), .cc2(\~ABL0 ));
SW0 switch1052 (.gate(\op-asl/rol ), .cc(net790));
SW0 switch1053 (.gate(notir2), .cc(\op-sty/cpy-mem ));
SW0 switch1054 (.gate(notir2), .cc(\op-T2-idx-x-xy ));
SW0 switch1055 (.gate(notir2), .cc(\op-T0-ldy-mem ));
SW0 switch1056 (.gate(notir2), .cc(\op-jmp ));
SW0 switch1057 (.gate(notir2), .cc(\op-T2-abs ));
SW0 switch1058 (.gate(notir2), .cc(\op-T3-jmp ));
SW0 switch1059 (.gate(notir2), .cc(\op-T0-bit ));
SW0 switch1060 (.gate(notir2), .cc(\op-T2-zp/zp-idx ));
SW0 switch1061 (.gate(notir2), .cc(\op-T0-jmp ));
SW0 switch1062 (.gate(notir2), .cc(\x-op-jmp ));
SW0 switch1063 (.gate(notir2), .cc(\op-T4-jmp ));
SW0 switch1064 (.gate(notir2), .cc(\op-T2-jmp-abs ));
SW0 switch1065 (.gate(notir2), .cc(\op-T+-bit ));
SW0 switch1066 (.gate(notir2), .cc(\op-T3-mem-zp-idx ));
SW0 switch1067 (.gate(notir2), .cc(\x-op-T0-bit ));
SW0 switch1068 (.gate(notir2), .cc(\op-T+-cpx/cpy-abs ));
SW0 switch1069 (.gate(notir2), .cc(\op-T3-mem-abs ));
SW0 switch1070 (.gate(notir2), .cc(\op-T2-mem-zp ));
SW0 switch1071 (.gate(cclk), .cc(dpc12_0ADD));
SW0 switch1072 (.gate(cclk), .cc(dpc11_SBADD));
SW0 switch1073 (.gate(cclk), .cc(dpc10_ADLADD));
SW0 switch1074 (.gate(cclk), .cc(dpc9_DBADD));
SW0 switch1075 (.gate(cclk), .cc(dpc8_nDBADD));
SW0 switch1076 (.gate(cclk), .cc(dpc7_SS));
SW0 switch1077 (.gate(cclk), .cc(dpc6_SBS));
SW0 switch1078 (.gate(dpc12_0ADD), .cc(alua0));
SW switch1079 (.gate(cp1), .cc1(\~TWOCYCLE ), .cc2(\~TWOCYCLE.phi1 ));
SW0 switch1080 (.gate(dpc12_0ADD), .cc(alua1));
SW0 switch1081 (.gate(dpc12_0ADD), .cc(alua4));
SW0 switch1082 (.gate(dpc12_0ADD), .cc(alua6));
SW0 switch1083 (.gate(dpc12_0ADD), .cc(alua5));
SW0 switch1084 (.gate(\x-op-jmp ), .cc(net510));
SW0 switch1085 (.gate(\x-op-jmp ), .cc(net134));
SW0 switch1086 (.gate(notalucin), .cc(net105));
SW0 switch1087 (.gate(notalucin), .cc(net942));
SW switch1088 (.gate(net37), .cc1(db2), .cc2(db2));
SW0 switch1089 (.gate(net37), .cc(db2));
SW0 switch1090 (.gate(net37), .cc(db2));
SW0 switch1091 (.gate(net37), .cc(db2));
SW0 switch1092 (.gate(net37), .cc(db2));
SW0 switch1093 (.gate(net37), .cc(db2));
SW0 switch1094 (.gate(net37), .cc(db2));
SW0 switch1095 (.gate(net37), .cc(db2));
SW0 switch1096 (.gate(net37), .cc(db2));
SW0 switch1097 (.gate(net8), .cc(net36));
SW0 switch1098 (.gate(net8), .cc(net150));
SW switch1099 (.gate(net570), .cc1(net1030), .cc2(DC78));
SW0 switch1100 (.gate(net1258), .cc(net591));
SW1 switch1101 (.gate(cclk), .cc(adl3));
SW0 switch1102 (.gate(\op-T4-ind-x ), .cc(net1649));
SW switch1103 (.gate(cclk), .cc1(net1724), .cc2(x6));
SW0 switch1104 (.gate(pipeUNK28), .cc(net1598));
SW0 switch1105 (.gate(net1238), .cc(dpc25_SBDB));
SW switch1106 (.gate(dpc17_SUMS), .cc1(\~(AxBxC)0 ), .cc2(\~aluresult0 ));
SW switch1107 (.gate(dpc17_SUMS), .cc1(\~(AxBxC)1 ), .cc2(\~aluresult1 ));
SW switch1108 (.gate(dpc17_SUMS), .cc1(\~(AxBxC)2 ), .cc2(\~aluresult2 ));
SW switch1109 (.gate(dpc17_SUMS), .cc1(\~(AxBxC)3 ), .cc2(\~aluresult3 ));
SW switch1110 (.gate(dpc17_SUMS), .cc1(\~(AxBxC)4 ), .cc2(\~aluresult4 ));
SW switch1111 (.gate(dpc17_SUMS), .cc1(\~(AxBxC)5 ), .cc2(\~aluresult5 ));
SW switch1112 (.gate(dpc17_SUMS), .cc1(\~aluresult6 ), .cc2(\~(AxBxC)6 ));
SW switch1113 (.gate(dpc17_SUMS), .cc1(\~aluresult7 ), .cc2(\~(AxBxC)7 ));
SW switch1114 (.gate(cp1), .cc1(net1376), .cc2(notdor2));
SW0 switch1115 (.gate(\x-op-T4-rti ), .cc(net327));
SW0 switch1116 (.gate(net988), .cc(AxB3));
SW switch1117 (.gate(cclk), .cc1(net34), .cc2(nots3));
SW1 switch1118 (.gate(cclk), .cc(sb3));
SW0 switch1119 (.gate(pipeUNK39), .cc(net2));
SW0 switch1120 (.gate(\~pclp5 ), .cc(pclp5));
SW switch1121 (.gate(cp1), .cc1(net1339), .cc2(net597));
SW0 switch1122 (.gate(net402), .cc(net834));
SW0 switch1123 (.gate(notx4), .cc(net436));
SW0 switch1124 (.gate(pd1), .cc(\pd1.clearIR ));
SW switch1125 (.gate(cclk), .cc1(net442), .cc2(net509));
SW0 switch1126 (.gate(noty0), .cc(net564));
SW0 switch1127 (.gate(notir7), .cc(\op-sty/cpy-mem ));
SW0 switch1128 (.gate(notir7), .cc(\op-T0-iny/dey ));
SW0 switch1129 (.gate(notir7), .cc(\x-op-T0-tya ));
SW0 switch1130 (.gate(notir7), .cc(\op-T0-cpy/iny ));
SW0 switch1131 (.gate(notir7), .cc(\op-xy ));
SW0 switch1132 (.gate(notir7), .cc(\x-op-T0-txa ));
SW0 switch1133 (.gate(notir7), .cc(\op-T0-dex ));
SW0 switch1134 (.gate(notir7), .cc(\op-T0-cpx/inx ));
SW0 switch1135 (.gate(notir7), .cc(\op-from-x ));
SW0 switch1136 (.gate(notir7), .cc(\op-T0-txs ));
SW0 switch1137 (.gate(notir7), .cc(\op-T0-ldx/tax/tsx ));
SW0 switch1138 (.gate(notir7), .cc(\op-T+-dex ));
SW0 switch1139 (.gate(notir7), .cc(\op-T+-inx ));
SW0 switch1140 (.gate(notir7), .cc(\op-T0-tsx ));
SW0 switch1141 (.gate(notir7), .cc(\op-T+-iny/dey ));
SW0 switch1142 (.gate(notir7), .cc(\op-T0-ldy-mem ));
SW0 switch1143 (.gate(notir7), .cc(\op-T0-tay/ldy-not-idx ));
SW0 switch1144 (.gate(notir7), .cc(\op-inc/nop ));
SW0 switch1145 (.gate(notir7), .cc(\op-T0-cpx/cpy/inx/iny ));
SW0 switch1146 (.gate(notir7), .cc(\op-T0-cmp ));
SW0 switch1147 (.gate(notir7), .cc(\op-T0-sbc ));
SW0 switch1148 (.gate(notir7), .cc(\op-T0-tya ));
SW0 switch1149 (.gate(notir7), .cc(\op-T0-txa ));
SW0 switch1150 (.gate(notir7), .cc(\op-T0-lda ));
SW0 switch1151 (.gate(notir7), .cc(\op-T0-tay ));
SW0 switch1152 (.gate(notir7), .cc(\op-T0-tax ));
SW0 switch1153 (.gate(notir7), .cc(\op-sta/cmp ));
SW0 switch1154 (.gate(notir7), .cc(\op-store ));
SW0 switch1155 (.gate(notir7), .cc(\op-T+-cmp ));
SW0 switch1156 (.gate(notir7), .cc(\op-T+-cpx/cpy-abs ));
SW0 switch1157 (.gate(notir7), .cc(\op-T+-cpx/cpy-imm/zp ));
SW0 switch1158 (.gate(notir7), .cc(\op-T0-cld/sed ));
SW0 switch1159 (.gate(notir7), .cc(\op-clv ));
SW switch1160 (.gate(dpc8_nDBADD), .cc1(alub0), .cc2(net624));
SW0 switch1161 (.gate(net236), .cc(net79));
SW0 switch1162 (.gate(C23), .cc(\~C23 ));
SW switch1163 (.gate(C23), .cc1(\~C34 ), .cc2(net924));
SW switch1164 (.gate(dpc8_nDBADD), .cc1(alub4), .cc2(net478));
SW switch1165 (.gate(dpc8_nDBADD), .cc1(alub2), .cc2(net458));
SW0 switch1166 (.gate(net811), .cc(net753));
SW0 switch1167 (.gate(net811), .cc(net753));
SW0 switch1168 (.gate(net519), .cc(net127));
SW1 switch1169 (.gate(net519), .cc(net135));
SW0 switch1170 (.gate(net1360), .cc(net1575));
SW0 switch1171 (.gate(\x-op-T+-adc/sbc ), .cc(\~op-set-C ));
SW0 switch1172 (.gate(\~A.B0 ), .cc(net1348));
SW switch1173 (.gate(net16), .cc1(net1703), .cc2(net468));
SW0 switch1174 (.gate(\op-T0-shift-right-a ), .cc(net366));
SW switch1175 (.gate(\~A.B4 ), .cc1(\~(AxB)4 ), .cc2(net1583));
SW0 switch1176 (.gate(\~ABL5 ), .cc(abl5));
SW0 switch1177 (.gate(net946), .cc(net384));
SW0 switch1178 (.gate(a7), .cc(net128));
SW0 switch1179 (.gate(net773), .cc(net275));
SW0 switch1180 (.gate(abl1), .cc(net66));
SW0 switch1181 (.gate(abl1), .cc(net842));
SW1 switch1182 (.gate(abl1), .cc(net1479));
SW switch1183 (.gate(cclk), .cc1(x1), .cc2(net1709));
SW0 switch1184 (.gate(\0/ADL1 ), .cc(adl1));
SW switch1185 (.gate(cp1), .cc1(net562), .cc2(net645));
SW0 switch1186 (.gate(net467), .cc(net1705));
SW switch1187 (.gate(net1392), .cc1(\~NMIP ), .cc2(net346));
SW0 switch1188 (.gate(net1392), .cc(net284));
SW0 switch1189 (.gate(net526), .cc(\~pclp0 ));
SW0 switch1190 (.gate(\op-T0-php/pha ), .cc(net1464));
SW0 switch1191 (.gate(\~C34 ), .cc(C34));
SW switch1192 (.gate(\~C34 ), .cc1(net1310), .cc2(C45));
SW0 switch1193 (.gate(\A+B7 ), .cc(net1617));
SW0 switch1194 (.gate(\~ABH3 ), .cc(abh3));
SW0 switch1195 (.gate(idb1), .cc(DBZ));
SW0 switch1196 (.gate(\PD-1xx000x0 ), .cc(\~TWOCYCLE ));
SW switch1197 (.gate(cclk), .cc1(pipeUNK37), .cc2(net944));
SW0 switch1198 (.gate(\op-T0-cpx/inx ), .cc(net1106));
SW switch1199 (.gate(cp1), .cc1(net1684), .cc2(notdor6));
SW0 switch1200 (.gate(\DA-AxB2 ), .cc(net388));
SW0 switch1201 (.gate(net1221), .cc(net1566));
SW0 switch1202 (.gate(net812), .cc(net1044));
SW switch1203 (.gate(cclk), .cc1(\~WR ), .cc2(\pipe~WR.phi2 ));
SW0 switch1204 (.gate(\op-T0-cmp ), .cc(net1560));
SW switch1205 (.gate(cp1), .cc1(net1375), .cc2(net95));
SW switch1206 (.gate(cp1), .cc1(net1089), .cc2(net1529));
SW switch1207 (.gate(net844), .cc1(net454), .cc2(net946));
SW switch1208 (.gate(dpc20_ADDSB06), .cc1(alu6), .cc2(sb6));
SW switch1209 (.gate(dpc20_ADDSB06), .cc1(alu5), .cc2(sb5));
SW switch1210 (.gate(dpc20_ADDSB06), .cc1(dasb4), .cc2(alu4));
SW switch1211 (.gate(dpc20_ADDSB06), .cc1(alu3), .cc2(sb3));
SW0 switch1212 (.gate(\op-T4-brk ), .cc(net1391));
SW0 switch1213 (.gate(\op-T4-brk ), .cc(\~WR ));
SW switch1214 (.gate(cclk), .cc1(\~pchp4 ), .cc2(net1657));
SW switch1215 (.gate(net553), .cc1(net511), .cc2(net845));
SW0 switch1216 (.gate(\notRdy0.phi1 ), .cc(net608));
SW0 switch1217 (.gate(adl0), .cc(net123));
SW0 switch1218 (.gate(alua4), .cc(net185));
SW0 switch1219 (.gate(alua4), .cc(\~(A+B)4 ));
SW0 switch1220 (.gate(net43), .cc(net21));
SW0 switch1221 (.gate(net1449), .cc(net944));
SW0 switch1222 (.gate(net1675), .cc(ir6));
SW switch1223 (.gate(net16), .cc1(net363), .cc2(net1091));
SW0 switch1224 (.gate(\op-T0-cpy/iny ), .cc(net1717));
SW0 switch1225 (.gate(net384), .cc(net885));
SW0 switch1226 (.gate(net384), .cc(net550));
SW switch1227 (.gate(cclk), .cc1(net176), .cc2(net598));
SW switch1228 (.gate(cclk), .cc1(net1592), .cc2(a7));
SW0 switch1229 (.gate(cclk), .cc(net891));
SW0 switch1230 (.gate(notir1), .cc(\op-xy ));
SW0 switch1231 (.gate(notir1), .cc(\x-op-T0-txa ));
SW0 switch1232 (.gate(notir1), .cc(\op-T0-dex ));
SW0 switch1233 (.gate(notir1), .cc(\op-from-x ));
SW0 switch1234 (.gate(notir1), .cc(\op-T0-txs ));
SW0 switch1235 (.gate(notir1), .cc(\op-T0-ldx/tax/tsx ));
SW0 switch1236 (.gate(notir1), .cc(\op-T+-dex ));
SW0 switch1237 (.gate(notir1), .cc(\op-T0-tsx ));
SW0 switch1238 (.gate(notir1), .cc(\op-ror ));
SW0 switch1239 (.gate(notir1), .cc(\op-inc/nop ));
SW0 switch1240 (.gate(notir1), .cc(\op-rol/ror ));
SW0 switch1241 (.gate(notir1), .cc(\op-shift ));
SW0 switch1242 (.gate(notir1), .cc(\op-T+-shift-a ));
SW0 switch1243 (.gate(notir1), .cc(\op-T0-txa ));
SW0 switch1244 (.gate(notir1), .cc(\op-T0-shift-a ));
SW0 switch1245 (.gate(notir1), .cc(\op-T0-tax ));
SW0 switch1246 (.gate(notir1), .cc(\op-T0-shift-right-a ));
SW0 switch1247 (.gate(notir1), .cc(\op-shift-right ));
SW0 switch1248 (.gate(notir1), .cc(\op-lsr/ror/dec/inc ));
SW0 switch1249 (.gate(notir1), .cc(\op-asl/rol ));
SW0 switch1250 (.gate(notir1), .cc(\op-T+-asl/rol-a ));
SW0 switch1251 (.gate(notRdy0), .cc(net191));
SW0 switch1252 (.gate(ONEBYTE), .cc(net1275));
SW0 switch1253 (.gate(net31), .cc(Pout0));
SW1 switch1254 (.gate(dor3), .cc(net42));
SW0 switch1255 (.gate(\op-ANDS ), .cc(\op-SUMS ));
SW1 switch1256 (.gate(net1140), .cc(ab9));
SW switch1257 (.gate(cclk), .cc1(RESP), .cc2(pipephi2Reset0x));
SW0 switch1258 (.gate(\~(A+B)5 ), .cc(\A+B5 ));
SW0 switch1259 (.gate(\~(A+B)5 ), .cc(AxB5));
SW0 switch1260 (.gate(net163), .cc(net1498));
SW0 switch1261 (.gate(net163), .cc(net903));
SW0 switch1262 (.gate(net1620), .cc(ir3));
SW switch1263 (.gate(cclk), .cc1(pipeUNK11), .cc2(net862));
SW switch1264 (.gate(cp1), .cc1(net1687), .cc2(notdor0));
SW switch1265 (.gate(cp1), .cc1(net299), .cc2(net1625));
SW switch1266 (.gate(cclk), .cc1(pipeUNK29), .cc2(net169));
SW0 switch1267 (.gate(pipeUNK26), .cc(net1714));
SW0 switch1268 (.gate(net1244), .cc(net1103));
SW0 switch1269 (.gate(net1433), .cc(net620));
SW switch1270 (.gate(cp1), .cc1(net254), .cc2(net1353));
SW switch1271 (.gate(cclk), .cc1(net340), .cc2(pipeUNK12));
SW switch1272 (.gate(\~A.B2 ), .cc1(net433), .cc2(C23));
SW switch1273 (.gate(net1446), .cc1(\short-circuit-branch-add ), .cc2(\~alucout ));
SW0 switch1274 (.gate(net1010), .cc(net311));
SW0 switch1275 (.gate(net1010), .cc(dpc35_PCHC));
SW0 switch1276 (.gate(net1047), .cc(dpc23_SBAC));
SW0 switch1277 (.gate(net796), .cc(net35));
SW switch1278 (.gate(net1262), .cc1(net1407), .cc2(net933));
SW switch1279 (.gate(cclk), .cc1(\~aluresult4 ), .cc2(notalu4));
SW0 switch1280 (.gate(\pd5.clearIR ), .cc(net928));
SW switch1281 (.gate(net284), .cc1(net891), .cc2(NMIP));
SW0 switch1282 (.gate(pch1), .cc(net1070));
SW0 switch1283 (.gate(notir4), .cc(\op-T3-ind-y ));
SW0 switch1284 (.gate(notir4), .cc(\op-T2-abs-y ));
SW0 switch1285 (.gate(notir4), .cc(\x-op-T0-tya ));
SW0 switch1286 (.gate(notir4), .cc(\op-T2-idx-x-xy ));
SW0 switch1287 (.gate(notir4), .cc(\op-T0-txs ));
SW0 switch1288 (.gate(notir4), .cc(\op-T0-tsx ));
SW0 switch1289 (.gate(notir4), .cc(\op-T4-ind-y ));
SW0 switch1290 (.gate(notir4), .cc(\op-T2-ind-y ));
SW0 switch1291 (.gate(notir4), .cc(\op-T3-abs-idx ));
SW0 switch1292 (.gate(notir4), .cc(\x-op-T3-ind-y ));
SW0 switch1293 (.gate(notir4), .cc(\op-T0-tya ));
SW0 switch1294 (.gate(notir4), .cc(\op-T4-abs-idx ));
SW0 switch1295 (.gate(notir4), .cc(\op-T5-ind-y ));
SW0 switch1296 (.gate(notir4), .cc(\op-branch-done ));
SW0 switch1297 (.gate(notir4), .cc(\op-T2-branch ));
SW0 switch1298 (.gate(notir4), .cc(\x-op-T4-ind-y ));
SW0 switch1299 (.gate(notir4), .cc(\x-op-T3-abs-idx ));
SW0 switch1300 (.gate(notir4), .cc(\op-T3-branch ));
SW0 switch1301 (.gate(notir4), .cc(\op-T0-cli/sei ));
SW0 switch1302 (.gate(notir4), .cc(\op-T0-clc/sec ));
SW0 switch1303 (.gate(notir4), .cc(\op-T3-mem-zp-idx ));
SW0 switch1304 (.gate(notir4), .cc(\op-T0-cld/sed ));
SW0 switch1305 (.gate(notir4), .cc(\op-T4-mem-abs-idx ));
SW0 switch1306 (.gate(notir4), .cc(\op-clv ));
SW0 switch1307 (.gate(adh2), .cc(net168));
SW switch1308 (.gate(dpc10_ADLADD), .cc1(adl2), .cc2(alub2));
SW switch1309 (.gate(cclk), .cc1(net889), .cc2(pipeUNK42));
SW0 switch1310 (.gate(idb1), .cc(net1474));
SW0 switch1311 (.gate(net1247), .cc(dpc30_ADHPCH));
SW0 switch1312 (.gate(net1247), .cc(dpc26_ACDB));
SW0 switch1313 (.gate(pipeUNK40), .cc(net1039));
SW0 switch1314 (.gate(net647), .cc(net939));
SW switch1315 (.gate(cclk), .cc1(\~ABL3 ), .cc2(net138));
SW0 switch1316 (.gate(pipephi2Reset0x), .cc(net717));
SW0 switch1317 (.gate(so), .cc(net1650));
SW0 switch1318 (.gate(net509), .cc(net1270));
SW0 switch1319 (.gate(net653), .cc(net390));
SW0 switch1320 (.gate(\op-T0-txa ), .cc(net1455));
SW0 switch1321 (.gate(net862), .cc(net1365));
SW1 switch1322 (.gate(net866), .cc(net9));
SW0 switch1323 (.gate(net1055), .cc(net1560));
SW0 switch1324 (.gate(net1038), .cc(net269));
SW0 switch1325 (.gate(\pd0.clearIR ), .cc(\PD-xxxx10x0 ));
SW0 switch1326 (.gate(\pd0.clearIR ), .cc(\PD-1xx000x0 ));
SW0 switch1327 (.gate(noty2), .cc(net1491));
SW0 switch1328 (.gate(net882), .cc(NMIL));
SW0 switch1329 (.gate(\dpc22_~DSA ), .cc(net306));
SW0 switch1330 (.gate(net1448), .cc(net1619));
SW switch1331 (.gate(cclk), .cc1(net831), .cc2(a5));
SW switch1332 (.gate(net1511), .cc1(net1598), .cc2(net262));
SW switch1333 (.gate(H1x1), .cc1(Pout1), .cc2(idb1));
SW0 switch1334 (.gate(net172), .cc(net1633));
SW1 switch1335 (.gate(net172), .cc(net210));
SW0 switch1336 (.gate(net1357), .cc(net678));
SW0 switch1337 (.gate(idb3), .cc(net1600));
SW switch1338 (.gate(dpc3_SBX), .cc1(x1), .cc2(sb1));
SW0 switch1339 (.gate(net1533), .cc(net964));
SW0 switch1340 (.gate(alu6), .cc(net149));
SW0 switch1341 (.gate(dpc12_0ADD), .cc(alua7));
SW0 switch1342 (.gate(net1715), .cc(net1399));
SW0 switch1343 (.gate(net1715), .cc(net1399));
SW1 switch1344 (.gate(net1715), .cc(net1105));
SW0 switch1345 (.gate(\op-T3-abs/idx/ind ), .cc(net726));
SW0 switch1346 (.gate(y4), .cc(noty4));
SW0 switch1347 (.gate(pcl1), .cc(net329));
SW0 switch1348 (.gate(net689), .cc(VEC0));
SW switch1349 (.gate(cclk), .cc1(net396), .cc2(net796));
SW switch1350 (.gate(cclk), .cc1(\~ABL0 ), .cc2(net1100));
SW0 switch1351 (.gate(pipeUNK13), .cc(net793));
SW0 switch1352 (.gate(net1380), .cc(net109));
SW0 switch1353 (.gate(nnT2BR), .cc(net405));
SW0 switch1354 (.gate(net1693), .cc(net1312));
SW0 switch1355 (.gate(\op-sty/cpy-mem ), .cc(net1604));
SW0 switch1356 (.gate(\op-sty/cpy-mem ), .cc(net1397));
SW0 switch1357 (.gate(net1247), .cc(dpc24_ACSB));
SW switch1359 (.gate(net269), .cc1(net1030), .cc2(DC78));
SW0 switch1360 (.gate(net603), .cc(\op-branch-done ));
SW switch1361 (.gate(alub6), .cc1(net1483), .cc2(\~A.B6 ));
SW0 switch1362 (.gate(alub6), .cc(\~(A+B)6 ));
SW0 switch1363 (.gate(net149), .cc(net970));
SW0 switch1364 (.gate(net149), .cc(net762));
SW0 switch1365 (.gate(idb4), .cc(net478));
SW0 switch1366 (.gate(\~(AxB1).C01 ), .cc(\~(AxBxC)1 ));
SW0 switch1367 (.gate(\op-push/pull ), .cc(\op-T2-abs-access ));
SW0 switch1368 (.gate(\op-push/pull ), .cc(\op-T3-abs/idx/ind ));
SW0 switch1369 (.gate(notidl0), .cc(idl0));
SW0 switch1370 (.gate(notidl0), .cc(idl0));
SW0 switch1371 (.gate(notidl0), .cc(idl0));
SW0 switch1372 (.gate(net1683), .cc(net966));
SW0 switch1373 (.gate(net441), .cc(dpc1_SBY));
SW0 switch1374 (.gate(net1109), .cc(net1649));
SW0 switch1375 (.gate(p1), .cc(net318));
SW switch1376 (.gate(net538), .cc1(net330), .cc2(net881));
SW0 switch1377 (.gate(net43), .cc(net1223));
SW0 switch1378 (.gate(net282), .cc(dpc6_SBS));
SW0 switch1379 (.gate(\~pchp5 ), .cc(pchp5));
SW0 switch1380 (.gate(net853), .cc(net1517));
SW0 switch1381 (.gate(AxB1), .cc(net1388));
SW0 switch1382 (.gate(AxB1), .cc(\~(AxB1).C01 ));
SW0 switch1383 (.gate(net876), .cc(net1584));
SW switch1384 (.gate(dpc37_PCLDB), .cc1(pclp6), .cc2(idb6));
SW0 switch1385 (.gate(net1356), .cc(net326));
SW0 switch1386 (.gate(\~A.B7 ), .cc(net637));
SW0 switch1387 (.gate(\~(A+B)2 ), .cc(\DA-AxB2 ));
SW0 switch1388 (.gate(notalu0), .cc(alu0));
SW0 switch1389 (.gate(dor6), .cc(net471));
SW0 switch1390 (.gate(dor6), .cc(net466));
SW switch1391 (.gate(cp1), .cc1(net1290), .cc2(net698));
SW switch1392 (.gate(cclk), .cc1(net111), .cc2(pd2));
SW switch1393 (.gate(cclk), .cc1(net62), .cc2(pd7));
SW switch1394 (.gate(cclk), .cc1(net374), .cc2(pd6));
SW0 switch1395 (.gate(IRQP), .cc(\~IRQP ));
SW0 switch1396 (.gate(IRQP), .cc(\~IRQP ));
SW0 switch1397 (.gate(notalu1), .cc(alu1));
SW0 switch1398 (.gate(\op-T2-branch ), .cc(net636));
SW switch1399 (.gate(\~TWOCYCLE.phi1 ), .cc1(net732), .cc2(net106));
SW0 switch1400 (.gate(db0), .cc(net93));
SW0 switch1401 (.gate(a2), .cc(net419));
SW0 switch1402 (.gate(ir7), .cc(notir7));
SW0 switch1403 (.gate(net1304), .cc(net1688));
SW0 switch1404 (.gate(nots3), .cc(net998));
SW0 switch1405 (.gate(notRdy0), .cc(net1145));
SW0 switch1406 (.gate(notRdy0), .cc(net604));
SW switch1407 (.gate(cp1), .cc1(net533), .cc2(net599));
SW0 switch1408 (.gate(nots1), .cc(net694));
SW0 switch1409 (.gate(net321), .cc(net849));
SW1 switch1410 (.gate(net321), .cc(dpc33_PCHDB));
SW0 switch1411 (.gate(\op-ANDS ), .cc(net384));
SW0 switch1412 (.gate(\op-ANDS ), .cc(net384));
SW0 switch1413 (.gate(net1377), .cc(net385));
SW0 switch1414 (.gate(net1177), .cc(net1614));
SW0 switch1415 (.gate(\op-rti/rts ), .cc(net300));
SW0 switch1416 (.gate(RnWstretched), .cc(net520));
SW0 switch1417 (.gate(RnWstretched), .cc(net520));
SW0 switch1418 (.gate(RnWstretched), .cc(net224));
SW0 switch1419 (.gate(notir0), .cc(\op-T3-ind-y ));
SW0 switch1420 (.gate(notir0), .cc(\op-T2-abs-y ));
SW0 switch1421 (.gate(notir0), .cc(\op-T2-ind-x ));
SW0 switch1422 (.gate(notir0), .cc(\op-T0-eor ));
SW0 switch1423 (.gate(notir0), .cc(\op-T0-ora ));
SW0 switch1424 (.gate(notir0), .cc(\op-T3-ind-x ));
SW0 switch1425 (.gate(notir0), .cc(\op-T4-ind-y ));
SW0 switch1426 (.gate(notir0), .cc(\op-T2-ind-y ));
SW0 switch1427 (.gate(notir0), .cc(\op-T4-ind-x ));
SW0 switch1428 (.gate(notir0), .cc(\x-op-T3-ind-y ));
SW0 switch1429 (.gate(notir0), .cc(\op-T0-cmp ));
SW0 switch1430 (.gate(notir0), .cc(\op-T0-sbc ));
SW0 switch1431 (.gate(notir0), .cc(\op-T0-adc/sbc ));
SW0 switch1432 (.gate(notir0), .cc(\op-T+-ora/and/eor/adc ));
SW0 switch1433 (.gate(notir0), .cc(\op-T+-adc/sbc ));
SW0 switch1434 (.gate(notir0), .cc(\op-T0-lda ));
SW0 switch1435 (.gate(notir0), .cc(\op-T0-acc ));
SW0 switch1436 (.gate(notir0), .cc(\op-T0-and ));
SW0 switch1437 (.gate(notir0), .cc(\op-T5-ind-y ));
SW0 switch1438 (.gate(notir0), .cc(\op-sta/cmp ));
SW0 switch1439 (.gate(notir0), .cc(\op-T2-ind ));
SW0 switch1440 (.gate(notir0), .cc(\op-T5-ind-x ));
SW0 switch1441 (.gate(notir0), .cc(\x-op-T4-ind-y ));
SW0 switch1442 (.gate(notir0), .cc(\x-op-T+-adc/sbc ));
SW0 switch1443 (.gate(notir0), .cc(\op-T+-cmp ));
SW0 switch1444 (.gate(notir0), .cc(\op-T5-mem-ind-idx ));
SW0 switch1446 (.gate(net759), .cc(net944));
SW switch1447 (.gate(fetch), .cc1(net1300), .cc2(net343));
SW0 switch1448 (.gate(\op-implied ), .cc(net664));
SW switch1449 (.gate(cp1), .cc1(IRQP), .cc2(net330));
SW0 switch1450 (.gate(RnWstretched), .cc(net612));
SW0 switch1451 (.gate(RnWstretched), .cc(net612));
SW switch1452 (.gate(cclk), .cc1(net14), .cc2(pipeUNK20));
SW switch1453 (.gate(cclk), .cc1(net586), .cc2(pipeUNK19));
SW0 switch1454 (.gate(t3), .cc(\op-T3-ind-y ));
SW0 switch1455 (.gate(t3), .cc(\op-T3-plp/pla ));
SW0 switch1456 (.gate(t3), .cc(\op-T3-stack/bit/jmp ));
SW0 switch1457 (.gate(t3), .cc(\op-T3-ind-x ));
SW0 switch1458 (.gate(t3), .cc(\op-T3-abs-idx ));
SW0 switch1459 (.gate(t3), .cc(\x-op-T3-ind-y ));
SW0 switch1460 (.gate(t3), .cc(\op-T3-jmp ));
SW0 switch1461 (.gate(t3), .cc(\op-T3-jsr ));
SW0 switch1462 (.gate(t3), .cc(\op-T3 ));
SW0 switch1463 (.gate(t3), .cc(\op-T3-abs/idx/ind ));
SW0 switch1464 (.gate(t3), .cc(\x-op-T3-abs-idx ));
SW0 switch1465 (.gate(t3), .cc(\op-T3-branch ));
SW0 switch1466 (.gate(t3), .cc(\x-op-T3-plp/pla ));
SW0 switch1467 (.gate(t3), .cc(\op-T3-mem-zp-idx ));
SW0 switch1468 (.gate(t3), .cc(\op-T3-mem-abs ));
SW switch1469 (.gate(net1682), .cc1(net613), .cc2(net150));
SW0 switch1470 (.gate(net91), .cc(net1256));
SW1 switch1471 (.gate(net91), .cc(dpc15_ANDS));
SW0 switch1472 (.gate(net339), .cc(net543));
SW0 switch1473 (.gate(net595), .cc(net239));
SW0 switch1474 (.gate(net595), .cc(net992));
SW0 switch1475 (.gate(net1247), .cc(dpc9_DBADD));
SW switch1476 (.gate(cclk), .cc1(net676), .cc2(\~ABH1 ));
SW1 switch1477 (.gate(net17), .cc(clock1));
SW0 switch1478 (.gate(net17), .cc(net646));
SW0 switch1479 (.gate(\op-T0-clc/sec ), .cc(net889));
SW0 switch1480 (.gate(\op-T0-plp ), .cc(net327));
SW switch1481 (.gate(\dpc41_DL/ADL ), .cc1(adl3), .cc2(net1661));
SW switch1482 (.gate(\dpc41_DL/ADL ), .cc1(adl4), .cc2(net1095));
SW switch1483 (.gate(\dpc41_DL/ADL ), .cc1(adl1), .cc2(net87));
SW switch1484 (.gate(\dpc41_DL/ADL ), .cc1(adl2), .cc2(net1424));
SW switch1485 (.gate(\dpc41_DL/ADL ), .cc1(adl0), .cc2(net719));
SW0 switch1486 (.gate(net320), .cc(net1322));
SW0 switch1487 (.gate(net320), .cc(net735));
SW0 switch1488 (.gate(RnWstretched), .cc(net471));
SW0 switch1489 (.gate(RnWstretched), .cc(net471));
SW0 switch1490 (.gate(\op-T4-abs-idx ), .cc(net595));
SW0 switch1491 (.gate(dor3), .cc(net643));
SW0 switch1492 (.gate(dor3), .cc(net1613));
SW switch1493 (.gate(cclk), .cc1(\pipe~VEC ), .cc2(\~VEC ));
SW0 switch1494 (.gate(\op-T0-brk/rti ), .cc(net256));
SW0 switch1495 (.gate(\A+B3 ), .cc(net924));
SW0 switch1496 (.gate(net1105), .cc(cp1));
SW0 switch1497 (.gate(net1105), .cc(cp1));
SW0 switch1498 (.gate(net1105), .cc(cp1));
SW0 switch1499 (.gate(net1105), .cc(cp1));
SW0 switch1500 (.gate(net1105), .cc(cp1));
SW0 switch1501 (.gate(net1488), .cc(net545));
SW0 switch1502 (.gate(net1488), .cc(net1547));
SW0 switch1503 (.gate(pipeVectorA2), .cc(net815));
SW0 switch1504 (.gate(net647), .cc(net570));
SW switch1505 (.gate(dpc0_YSB), .cc1(net1491), .cc2(sb2));
SW0 switch1506 (.gate(net470), .cc(net467));
SW switch1507 (.gate(cclk), .cc1(net146), .cc2(a0));
SW switch1508 (.gate(dpc0_YSB), .cc1(sb3), .cc2(net1531));
SW0 switch1509 (.gate(net885), .cc(net513));
SW0 switch1510 (.gate(RnWstretched), .cc(net37));
SW0 switch1511 (.gate(RnWstretched), .cc(net37));
SW switch1512 (.gate(alub3), .cc1(\~A.B3 ), .cc2(net313));
SW0 switch1513 (.gate(alub3), .cc(\~(A+B)3 ));
SW0 switch1514 (.gate(net288), .cc(net798));
SW1 switch1515 (.gate(net288), .cc(net794));
SW1 switch1516 (.gate(abh0), .cc(net826));
SW0 switch1517 (.gate(net43), .cc(net625));
SW0 switch1518 (.gate(s3), .cc(net34));
SW0 switch1519 (.gate(\~pchp6 ), .cc(pchp6));
SW0 switch1520 (.gate(net1677), .cc(net475));
SW1 switch1521 (.gate(net1677), .cc(net999));
SW switch1522 (.gate(cclk), .cc1(net865), .cc2(net958));
SW switch1523 (.gate(dpc3_SBX), .cc1(dasb4), .cc2(x4));
SW switch1524 (.gate(dpc3_SBX), .cc1(x3), .cc2(sb3));
SW switch1525 (.gate(dpc3_SBX), .cc1(x2), .cc2(sb2));
SW0 switch1526 (.gate(net582), .cc(net1067));
SW1 switch1527 (.gate(net582), .cc(\ADH/ABH ));
SW switch1528 (.gate(dpc3_SBX), .cc1(sb6), .cc2(x6));
SW switch1529 (.gate(dpc3_SBX), .cc1(x5), .cc2(sb5));
SW0 switch1530 (.gate(net1629), .cc(dasb5));
SW0 switch1531 (.gate(\~ABL2 ), .cc(abl2));
SW0 switch1532 (.gate(net71), .cc(dpc7_SS));
SW switch1533 (.gate(dpc3_SBX), .cc1(x7), .cc2(sb7));
SW0 switch1534 (.gate(a5), .cc(net1719));
SW0 switch1535 (.gate(\op-T3-ind-y ), .cc(net1717));
SW1 switch1536 (.gate(net520), .cc(db2));
SW1 switch1537 (.gate(net520), .cc(db2));
SW0 switch1538 (.gate(pipeUNK42), .cc(net253));
SW0 switch1539 (.gate(net1552), .cc(dpc14_SRS));
SW0 switch1540 (.gate(idb4), .cc(net797));
SW0 switch1541 (.gate(net644), .cc(net678));
SW0 switch1542 (.gate(net975), .cc(net854));
SW0 switch1543 (.gate(\~(A+B)6 ), .cc(\A+B6 ));
SW0 switch1544 (.gate(\~(A+B)6 ), .cc(C67));
SW switch1545 (.gate(net1205), .cc1(net1454), .cc2(dasb7));
SW0 switch1546 (.gate(net1205), .cc(net260));
SW switch1547 (.gate(cclk), .cc1(\op-EORS ), .cc2(net982));
SW1 switch1548 (.gate(cclk), .cc(sb7));
SW switch1549 (.gate(cclk), .cc1(\op-ORS ), .cc2(net88));
SW switch1550 (.gate(net1386), .cc1(net484), .cc2(net914));
SW0 switch1551 (.gate(net31), .cc(net307));
SW0 switch1552 (.gate(sb2), .cc(net1580));
SW0 switch1553 (.gate(sb2), .cc(net1580));
SW0 switch1554 (.gate(net86), .cc(ab4));
SW0 switch1555 (.gate(net86), .cc(ab4));
SW0 switch1556 (.gate(net86), .cc(ab4));
SW0 switch1557 (.gate(net86), .cc(ab4));
SW switch1558 (.gate(cp1), .cc1(net1624), .cc2(notRdy0));
SW0 switch1559 (.gate(\op-T0-tay/ldy-not-idx ), .cc(net616));
SW0 switch1560 (.gate(\A+B6 ), .cc(net482));
SW0 switch1561 (.gate(net210), .cc(ab5));
SW0 switch1562 (.gate(net210), .cc(ab5));
SW0 switch1563 (.gate(net210), .cc(ab5));
SW0 switch1564 (.gate(net210), .cc(ab5));
SW0 switch1565 (.gate(pipeUNK20), .cc(net959));
SW0 switch1566 (.gate(net128), .cc(net1592));
SW0 switch1567 (.gate(RnWstretched), .cc(net42));
SW0 switch1568 (.gate(RnWstretched), .cc(net42));
SW0 switch1569 (.gate(RnWstretched), .cc(net1613));
SW0 switch1570 (.gate(alucin), .cc(notalucin));
SW switch1571 (.gate(cclk), .cc1(net658), .cc2(y4));
SW0 switch1572 (.gate(net673), .cc(net1304));
SW0 switch1573 (.gate(net15), .cc(\~pclp4 ));
SW switch1574 (.gate(cp1), .cc1(net1514), .cc2(net880));
SW0 switch1575 (.gate(net708), .cc(dpc11_SBADD));
SW switch1576 (.gate(cclk), .cc1(y3), .cc2(net1531));
SW switch1577 (.gate(net480), .cc1(net202), .cc2(net629));
SW switch1578 (.gate(cp1), .cc1(net472), .cc2(net1606));
SW switch1579 (.gate(cclk), .cc1(pipeUNK05), .cc2(net90));
SW0 switch1580 (.gate(pipedpc28), .cc(dpc28_0ADH0));
SW0 switch1581 (.gate(net1154), .cc(net1380));
SW0 switch1582 (.gate(\op-T3-mem-zp-idx ), .cc(net347));
SW switch1583 (.gate(cclk), .cc1(\~notRdy0.delay ), .cc2(net608));
SW0 switch1584 (.gate(RnWstretched), .cc(net373));
SW0 switch1585 (.gate(RnWstretched), .cc(net373));
SW0 switch1586 (.gate(RnWstretched), .cc(net1720));
SW1 switch1587 (.gate(cclk), .cc(dasb0));
SW switch1588 (.gate(cclk), .cc1(\~aluresult6 ), .cc2(notalu6));
SW0 switch1589 (.gate(net409), .cc(\PD-xxx010x1 ));
SW switch1590 (.gate(dpc14_SRS), .cc1(\~A.B1 ), .cc2(\~aluresult0 ));
SW switch1591 (.gate(dpc14_SRS), .cc1(\~aluresult1 ), .cc2(\~A.B2 ));
SW switch1592 (.gate(dpc14_SRS), .cc1(\~A.B3 ), .cc2(\~aluresult2 ));
SW switch1593 (.gate(dpc14_SRS), .cc1(\~aluresult3 ), .cc2(\~A.B4 ));
SW switch1594 (.gate(dpc14_SRS), .cc1(\~aluresult4 ), .cc2(\~A.B5 ));
SW switch1595 (.gate(dpc14_SRS), .cc1(\~aluresult5 ), .cc2(\~A.B6 ));
SW switch1596 (.gate(dpc14_SRS), .cc1(\~aluresult6 ), .cc2(\~A.B7 ));
SW switch1597 (.gate(cclk), .cc1(net469), .cc2(net875));
SW0 switch1598 (.gate(\op-T+-inx ), .cc(net844));
SW switch1599 (.gate(dpc1_SBY), .cc1(y2), .cc2(sb2));
SW switch1600 (.gate(net613), .cc1(net1656), .cc2(dasb2));
SW0 switch1601 (.gate(net613), .cc(net1159));
SW1 switch1602 (.gate(cclk), .cc(idb7));
SW switch1603 (.gate(cclk), .cc1(VEC1), .cc2(net1452));
SW switch1604 (.gate(cclk), .cc1(\C78.phi2 ), .cc2(alurawcout));
SW0 switch1605 (.gate(net572), .cc(net1517));
SW switch1606 (.gate(\A+B0 ), .cc1(net1348), .cc2(\~(AxB)0 ));
SW0 switch1607 (.gate(net139), .cc(net169));
SW0 switch1608 (.gate(net334), .cc(Pout2));
SW0 switch1609 (.gate(RnWstretched), .cc(net643));
SW0 switch1610 (.gate(RnWstretched), .cc(net643));
SW0 switch1611 (.gate(notRdy0), .cc(net46));
SW0 switch1612 (.gate(net1137), .cc(\short-circuit-idx-add ));
SW0 switch1613 (.gate(\C78.phi2 ), .cc(notalucout));
SW0 switch1614 (.gate(\~(AxB3).C23 ), .cc(\~(AxBxC)3 ));
SW switch1615 (.gate(cclk), .cc1(net436), .cc2(x4));
SW switch1616 (.gate(cclk), .cc1(net896), .cc2(notidl3));
SW0 switch1617 (.gate(net1716), .cc(net180));
SW0 switch1618 (.gate(db7), .cc(net588));
SW0 switch1619 (.gate(net1045), .cc(Pout7));
SW switch1620 (.gate(cclk), .cc1(pipeUNK26), .cc2(net132));
SW switch1621 (.gate(cclk), .cc1(net1254), .cc2(\~ABL6 ));
SW0 switch1622 (.gate(net550), .cc(net1347));
SW switch1623 (.gate(net790), .cc1(net1137), .cc2(net816));
SW switch1624 (.gate(cclk), .cc1(\~aluresult1 ), .cc2(notalu1));
SW switch1625 (.gate(\ADL/ABL ), .cc1(\~ABL3 ), .cc2(net864));
SW0 switch1626 (.gate(db5), .cc(net1588));
SW0 switch1627 (.gate(net747), .cc(net1417));
SW0 switch1628 (.gate(\pd6.clearIR ), .cc(net1309));
SW0 switch1629 (.gate(\~op-branch-bit7 ), .cc(net201));
SW0 switch1630 (.gate(RnWstretched), .cc(net798));
SW0 switch1631 (.gate(RnWstretched), .cc(net798));
SW0 switch1632 (.gate(RnWstretched), .cc(net288));
SW0 switch1633 (.gate(cclk), .cc(net525));
SW0 switch1634 (.gate(cclk), .cc(net628));
SW0 switch1635 (.gate(net1111), .cc(net1470));
SW0 switch1636 (.gate(net1111), .cc(net1614));
SW0 switch1637 (.gate(alua3), .cc(net313));
SW0 switch1638 (.gate(alua3), .cc(\~(A+B)3 ));
SW0 switch1639 (.gate(net956), .cc(dpc12_0ADD));
SW0 switch1640 (.gate(notx3), .cc(net242));
SW switch1641 (.gate(dpc1_SBY), .cc1(y1), .cc2(sb1));
SW switch1642 (.gate(net440), .cc1(net137), .cc2(net504));
SW0 switch1643 (.gate(\brk-done ), .cc(net1649));
SW0 switch1644 (.gate(\brk-done ), .cc(net300));
SW0 switch1645 (.gate(net90), .cc(net1433));
SW0 switch1646 (.gate(\op-T3 ), .cc(net256));
SW switch1647 (.gate(alub4), .cc1(\~A.B4 ), .cc2(net185));
SW0 switch1648 (.gate(alub4), .cc(\~(A+B)4 ));
SW0 switch1649 (.gate(net1258), .cc(\~WR ));
SW0 switch1650 (.gate(notx0), .cc(net1169));
SW0 switch1651 (.gate(net95), .cc(net531));
SW switch1652 (.gate(cclk), .cc1(net31), .cc2(pipeUNK16));
SW switch1653 (.gate(cp1), .cc1(net1368), .cc2(net1149));
SW0 switch1654 (.gate(dor5), .cc(net612));
SW0 switch1655 (.gate(dor5), .cc(net1720));
SW0 switch1656 (.gate(net126), .cc(\~pchp1 ));
SW0 switch1657 (.gate(\op-T2-php ), .cc(net1391));
SW0 switch1658 (.gate(AxB3), .cc(net1610));
SW0 switch1659 (.gate(\~(AxB7).C67 ), .cc(\~(AxBxC)7 ));
SW0 switch1660 (.gate(net43), .cc(net476));
SW0 switch1661 (.gate(net453), .cc(net1213));
SW0 switch1662 (.gate(net1371), .cc(net620));
SW0 switch1663 (.gate(Pout3), .cc(net51));
SW0 switch1664 (.gate(p2), .cc(net334));
SW0 switch1665 (.gate(net1002), .cc(net605));
SW0 switch1666 (.gate(net1002), .cc(net605));
SW0 switch1667 (.gate(net1477), .cc(net1541));
SW0 switch1668 (.gate(\op-T3-ind-x ), .cc(net1107));
SW0 switch1669 (.gate(\op-T3-ind-x ), .cc(net604));
SW0 switch1671 (.gate(net646), .cc(net272));
SW0 switch1672 (.gate(\~op-branch-bit7 ), .cc(net1293));
SW0 switch1673 (.gate(\op-T0-pla ), .cc(net1455));
SW0 switch1674 (.gate(net800), .cc(dpc26_ACDB));
SW0 switch1675 (.gate(net1247), .cc(dpc31_PCHPCH));
SW switch1676 (.gate(\dpc41_DL/ADL ), .cc1(adl6), .cc2(net1014));
SW switch1677 (.gate(\dpc41_DL/ADL ), .cc1(adl5), .cc2(net1387));
SW switch1678 (.gate(cclk), .cc1(net1037), .cc2(net266));
SW1 switch1679 (.gate(net42), .cc(db3));
SW1 switch1680 (.gate(net42), .cc(db3));
SW0 switch1681 (.gate(s4), .cc(net973));
SW0 switch1682 (.gate(net1471), .cc(Pout4));
SW switch1683 (.gate(cclk), .cc1(net1586), .cc2(net621));
SW switch1684 (.gate(cp1), .cc1(net577), .cc2(net1046));
SW0 switch1685 (.gate(net476), .cc(net956));
SW1 switch1686 (.gate(net476), .cc(dpc12_0ADD));
SW0 switch1687 (.gate(\op-xy ), .cc(net1244));
SW0 switch1688 (.gate(\op-xy ), .cc(net1351));
SW0 switch1689 (.gate(idb5), .cc(net961));
SW switch1690 (.gate(cp1), .cc1(net1093), .cc2(net226));
SW0 switch1691 (.gate(\op-T0-txs ), .cc(net1358));
SW0 switch1692 (.gate(net671), .cc(net14));
SW0 switch1693 (.gate(net1124), .cc(net1662));
SW0 switch1694 (.gate(net1269), .cc(net1401));
SW0 switch1695 (.gate(net1269), .cc(net1249));
SW switch1696 (.gate(\ADH/ABH ), .cc1(\~ABH4 ), .cc2(net1451));
SW0 switch1697 (.gate(net226), .cc(net1593));
SW0 switch1698 (.gate(net543), .cc(net196));
SW1 switch1699 (.gate(net543), .cc(dpc5_SADL));
SW0 switch1700 (.gate(\~op-T3-branch ), .cc(net236));
SW1 switch1701 (.gate(net475), .cc(ab12));
SW0 switch1702 (.gate(INTG), .cc(D1x1));
SW switch1703 (.gate(cp1), .cc1(D1x1), .cc2(net1472));
SW switch1704 (.gate(cp1), .cc1(net1275), .cc2(net1581));
SW0 switch1705 (.gate(ir1), .cc(net1133));
SW0 switch1706 (.gate(ir1), .cc(notir1));
SW switch1707 (.gate(\ADH/ABH ), .cc1(\~ABH5 ), .cc2(net1353));
SW0 switch1708 (.gate(\op-T2-pha ), .cc(net1037));
SW0 switch1709 (.gate(net1399), .cc(net1105));
SW0 switch1710 (.gate(net319), .cc(net972));
SW0 switch1711 (.gate(net936), .cc(AxB1));
SW1 switch1712 (.gate(net1325), .cc(db0));
SW1 switch1713 (.gate(net1325), .cc(db0));
SW0 switch1714 (.gate(net43), .cc(net611));
SW0 switch1715 (.gate(\op-T0-txs ), .cc(net1106));
SW switch1716 (.gate(cp1), .cc1(net50), .cc2(INTG));
SW0 switch1717 (.gate(net600), .cc(net36));
SW0 switch1718 (.gate(\op-branch-done ), .cc(\~op-branch-done ));
SW switch1719 (.gate(cp1), .cc1(net1636), .cc2(net935));
SW0 switch1720 (.gate(notir5), .cc(net503));
SW switch1721 (.gate(dpc5_SADL), .cc1(adl5), .cc2(net280));
SW switch1722 (.gate(dpc5_SADL), .cc1(adl4), .cc2(net3));
SW switch1723 (.gate(dpc5_SADL), .cc1(adl3), .cc2(net998));
SW switch1724 (.gate(dpc5_SADL), .cc1(adl2), .cc2(net1389));
SW0 switch1725 (.gate(net1408), .cc(net1004));
SW0 switch1726 (.gate(net1662), .cc(net553));
SW switch1727 (.gate(dpc5_SADL), .cc1(net721), .cc2(adl7));
SW0 switch1728 (.gate(net862), .cc(net1347));
SW0 switch1729 (.gate(\~ABL1 ), .cc(abl1));
SW switch1730 (.gate(net236), .cc1(net182), .cc2(net1151));
SW0 switch1731 (.gate(\~pchp3 ), .cc(pchp3));
SW switch1732 (.gate(cp1), .cc1(net1528), .cc2(net1215));
SW switch1733 (.gate(cp1), .cc1(net1161), .cc2(net109));
SW switch1734 (.gate(net1401), .cc1(\branch-back ), .cc2(net1198));
SW0 switch1735 (.gate(notidl7), .cc(idl7));
SW0 switch1736 (.gate(notidl7), .cc(idl7));
SW0 switch1737 (.gate(notidl7), .cc(idl7));
SW0 switch1738 (.gate(\notRdy0.delay ), .cc(net19));
SW1 switch1739 (.gate(cclk), .cc(sb1));
SW switch1740 (.gate(cclk), .cc1(net182), .cc2(net265));
SW switch1741 (.gate(cclk), .cc1(net897), .cc2(net1211));
SW0 switch1742 (.gate(\op-T5-rti/rts ), .cc(net368));
SW0 switch1743 (.gate(notalucin), .cc(net1354));
SW0 switch1744 (.gate(net1214), .cc(fetch));
SW0 switch1745 (.gate(net966), .cc(net1635));
SW1 switch1746 (.gate(net966), .cc(dpc29_0ADH17));
SW0 switch1747 (.gate(\~notRdy0.delay ), .cc(\notRdy0.delay ));
SW0 switch1748 (.gate(net1596), .cc(net1271));
SW1 switch1749 (.gate(net1596), .cc(dpc27_SBADH));
SW1 switch1750 (.gate(cclk), .cc(adl2));
SW switch1751 (.gate(cclk), .cc1(net1402), .cc2(\~pchp2 ));
SW switch1752 (.gate(cp1), .cc1(net1014), .cc2(idl6));
SW switch1753 (.gate(net1600), .cc1(net1546), .cc2(net1495));
SW0 switch1754 (.gate(net31), .cc(net1044));
SW0 switch1755 (.gate(net905), .cc(net979));
SW0 switch1756 (.gate(net1533), .cc(clock2));
SW1 switch1757 (.gate(net373), .cc(db5));
SW1 switch1758 (.gate(net373), .cc(db5));
SW0 switch1759 (.gate(net1175), .cc(net267));
SW1 switch1760 (.gate(cclk), .cc(idb2));
SW0 switch1761 (.gate(net597), .cc(net882));
SW0 switch1762 (.gate(net761), .cc(net1056));
SW switch1763 (.gate(C34), .cc1(net695), .cc2(net619));
SW0 switch1764 (.gate(C34), .cc(net1179));
SW switch1765 (.gate(cclk), .cc1(net674), .cc2(net745));
SW switch1766 (.gate(cclk), .cc1(net1130), .cc2(net512));
SW switch1767 (.gate(cclk), .cc1(\~pclp1 ), .cc2(net1099));
SW0 switch1768 (.gate(AxB7), .cc(net269));
SW0 switch1769 (.gate(RnWstretched), .cc(net298));
SW0 switch1770 (.gate(RnWstretched), .cc(net298));
SW0 switch1771 (.gate(RnWstretched), .cc(net23));
SW0 switch1772 (.gate(net600), .cc(net1279));
SW0 switch1773 (.gate(net161), .cc(net969));
SW1 switch1774 (.gate(net161), .cc(dpc0_YSB));
SW0 switch1775 (.gate(net641), .cc(net715));
SW0 switch1776 (.gate(net641), .cc(dpc34_PCLC));
SW0 switch1777 (.gate(net1247), .cc(dpc7_SS));
SW0 switch1778 (.gate(\op-T4-brk/jsr ), .cc(net604));
SW switch1779 (.gate(dpc1_SBY), .cc1(y5), .cc2(sb5));
SW0 switch1780 (.gate(pipeUNK15), .cc(H1x1));
SW0 switch1781 (.gate(net1043), .cc(dpc40_ADLPCL));
SW switch1782 (.gate(dpc1_SBY), .cc1(y7), .cc2(sb7));
SW0 switch1783 (.gate(net1218), .cc(net1257));
SW0 switch1784 (.gate(pd3), .cc(\pd3.clearIR ));
SW0 switch1785 (.gate(db4), .cc(net490));
SW switch1786 (.gate(net344), .cc1(net1073), .cc2(net557));
SW1 switch1787 (.gate(net826), .cc(ab8));
SW switch1788 (.gate(net344), .cc1(net20), .cc2(net585));
SW0 switch1789 (.gate(net344), .cc(net1316));
SW switch1790 (.gate(cclk), .cc1(pipeUNK27), .cc2(\op-SRS ));
SW0 switch1791 (.gate(notRdy0), .cc(VEC0));
SW0 switch1792 (.gate(net1501), .cc(db7));
SW0 switch1793 (.gate(net1501), .cc(db7));
SW0 switch1794 (.gate(net1501), .cc(db7));
SW0 switch1795 (.gate(net1501), .cc(db7));
SW switch1796 (.gate(cclk), .cc1(net1049), .cc2(net160));
SW0 switch1797 (.gate(\~A.B5 ), .cc(net647));
SW0 switch1798 (.gate(net1149), .cc(\~NMIG ));
SW0 switch1799 (.gate(net1565), .cc(net1218));
SW0 switch1800 (.gate(net1565), .cc(net1218));
SW switch1801 (.gate(cp1), .cc1(notRdy0), .cc2(net1276));
SW switch1802 (.gate(cclk), .cc1(pipeUNK35), .cc2(net501));
SW0 switch1803 (.gate(t2), .cc(\op-T2-abs-y ));
SW0 switch1804 (.gate(t2), .cc(\op-T2-idx-x-xy ));
SW0 switch1805 (.gate(t2), .cc(\op-T2-ind-x ));
SW0 switch1806 (.gate(t2), .cc(\op-T2 ));
SW0 switch1807 (.gate(t2), .cc(\op-T2-abs ));
SW0 switch1808 (.gate(t2), .cc(\op-T2-ADL/ADD ));
SW0 switch1809 (.gate(t2), .cc(\op-T2-stack ));
SW0 switch1810 (.gate(t2), .cc(\op-T2-ind-y ));
SW0 switch1811 (.gate(t2), .cc(\op-T2-jsr ));
SW0 switch1812 (.gate(t2), .cc(\op-T2-stack-access ));
SW0 switch1813 (.gate(t2), .cc(\op-T2-pha ));
SW0 switch1814 (.gate(t2), .cc(\op-T2-brk ));
SW0 switch1815 (.gate(t2), .cc(\op-T2-branch ));
SW0 switch1816 (.gate(t2), .cc(\op-T2-zp/zp-idx ));
SW0 switch1817 (.gate(t2), .cc(\op-T2-ind ));
SW0 switch1818 (.gate(t2), .cc(\op-T2-abs-access ));
SW0 switch1819 (.gate(t2), .cc(\op-T2-php ));
SW0 switch1820 (.gate(t2), .cc(\op-T2-php/pha ));
SW0 switch1821 (.gate(t2), .cc(\op-T2-jmp-abs ));
SW0 switch1822 (.gate(t2), .cc(\op-T2-mem-zp ));
SW switch1823 (.gate(cp1), .cc1(net1360), .cc2(net1091));
SW0 switch1824 (.gate(\op-T2-ind-x ), .cc(net1106));
SW0 switch1825 (.gate(net1679), .cc(net1262));
SW switch1826 (.gate(cclk), .cc1(pipeUNK41), .cc2(net504));
SW switch1827 (.gate(cclk), .cc1(\op-ANDS ), .cc2(net1574));
SW0 switch1828 (.gate(y7), .cc(noty7));
SW switch1829 (.gate(cclk), .cc1(net119), .cc2(notir1));
SW0 switch1830 (.gate(ir0), .cc(\op-implied ));
SW switch1831 (.gate(fetch), .cc1(net237), .cc2(net119));
SW switch1832 (.gate(fetch), .cc1(net724), .cc2(net310));
SW switch1833 (.gate(cp1), .cc1(notRdy0), .cc2(\notRdy0.phi1 ));
SW0 switch1834 (.gate(net503), .cc(net270));
SW0 switch1835 (.gate(idb6), .cc(net1684));
SW0 switch1836 (.gate(\op-T5-rts ), .cc(net256));
SW switch1837 (.gate(net335), .cc1(net508), .cc2(net1303));
SW0 switch1838 (.gate(pd6), .cc(\pd6.clearIR ));
SW switch1839 (.gate(alub2), .cc1(\~A.B2 ), .cc2(net452));
SW0 switch1840 (.gate(alub2), .cc(\~(A+B)2 ));
SW switch1841 (.gate(dpc23_SBAC), .cc1(dasb0), .cc2(a0));
SW switch1842 (.gate(dpc23_SBAC), .cc1(dasb1), .cc2(a1));
SW switch1843 (.gate(dpc23_SBAC), .cc1(a2), .cc2(dasb2));
SW switch1844 (.gate(dpc23_SBAC), .cc1(dasb3), .cc2(a3));
SW switch1845 (.gate(dpc23_SBAC), .cc1(dasb4), .cc2(a4));
SW switch1846 (.gate(dpc23_SBAC), .cc1(dasb5), .cc2(a5));
SW switch1847 (.gate(dpc23_SBAC), .cc1(dasb6), .cc2(a6));
SW switch1848 (.gate(dpc23_SBAC), .cc1(dasb7), .cc2(a7));
SW0 switch1849 (.gate(net251), .cc(net1028));
SW0 switch1850 (.gate(net251), .cc(RnWstretched));
SW0 switch1851 (.gate(net251), .cc(RnWstretched));
SW0 switch1852 (.gate(net251), .cc(RnWstretched));
SW0 switch1853 (.gate(net251), .cc(RnWstretched));
SW0 switch1854 (.gate(\~op-T3-branch ), .cc(net19));
SW switch1855 (.gate(dpc25_SBDB), .cc1(dasb0), .cc2(idb0));
SW switch1856 (.gate(dpc25_SBDB), .cc1(sb1), .cc2(idb1));
SW switch1857 (.gate(dpc25_SBDB), .cc1(idb2), .cc2(sb2));
SW switch1858 (.gate(dpc25_SBDB), .cc1(sb3), .cc2(idb3));
SW switch1859 (.gate(dpc25_SBDB), .cc1(idb4), .cc2(dasb4));
SW switch1860 (.gate(dpc25_SBDB), .cc1(idb5), .cc2(sb5));
SW switch1861 (.gate(dpc25_SBDB), .cc1(idb6), .cc2(sb6));
SW switch1862 (.gate(dpc25_SBDB), .cc1(sb7), .cc2(idb7));
SW switch1863 (.gate(cclk), .cc1(net1065), .cc2(net1124));
SW0 switch1864 (.gate(\~C45 ), .cc(\DA-C45 ));
SW0 switch1865 (.gate(net1194), .cc(Pout3));
SW0 switch1866 (.gate(pipeUNK33), .cc(net1178));
SW switch1867 (.gate(cclk), .cc1(net824), .cc2(net398));
SW0 switch1868 (.gate(VEC0), .cc(net728));
SW switch1869 (.gate(net388), .cc1(net972), .cc2(DC34));
SW0 switch1870 (.gate(\~ABL3 ), .cc(abl3));
SW0 switch1871 (.gate(cclk), .cc(net742));
SW0 switch1872 (.gate(net616), .cc(net454));
SW0 switch1873 (.gate(\op-T0-cld/sed ), .cc(net774));
SW0 switch1874 (.gate(net390), .cc(net1258));
SW0 switch1875 (.gate(notdor6), .cc(dor6));
SW switch1876 (.gate(\dpc41_DL/ADL ), .cc1(net1147), .cc2(adl7));
SW0 switch1877 (.gate(net620), .cc(net922));
SW0 switch1878 (.gate(net620), .cc(net1115));
SW0 switch1879 (.gate(net1295), .cc(net1238));
SW1 switch1880 (.gate(net1295), .cc(dpc25_SBDB));
SW switch1881 (.gate(cclk), .cc1(net1209), .cc2(net663));
SW switch1882 (.gate(cp1), .cc1(net1181), .cc2(net69));
SW switch1883 (.gate(cclk), .cc1(\~ABL7 ), .cc2(net171));
SW0 switch1884 (.gate(net1247), .cc(dpc10_ADLADD));
SW0 switch1885 (.gate(\op-T+-cpx/cpy-imm/zp ), .cc(\~op-set-C ));
SW0 switch1886 (.gate(net799), .cc(net1339));
SW0 switch1887 (.gate(net643), .cc(db3));
SW0 switch1888 (.gate(net643), .cc(db3));
SW0 switch1889 (.gate(net643), .cc(db3));
SW0 switch1890 (.gate(net643), .cc(db3));
SW0 switch1891 (.gate(net643), .cc(db3));
SW0 switch1892 (.gate(net643), .cc(db3));
SW0 switch1893 (.gate(net643), .cc(db3));
SW1 switch1894 (.gate(net102), .cc(rw));
SW1 switch1895 (.gate(net102), .cc(rw));
SW1 switch1896 (.gate(net102), .cc(rw));
SW1 switch1897 (.gate(net102), .cc(rw));
SW1 switch1898 (.gate(net102), .cc(rw));
SW1 switch1899 (.gate(net102), .cc(rw));
SW1 switch1900 (.gate(net102), .cc(rw));
SW0 switch1901 (.gate(C67), .cc(\~C67 ));
SW switch1902 (.gate(C67), .cc1(\~C78 ), .cc2(net1617));
SW0 switch1903 (.gate(net1083), .cc(\PD-xxx010x1 ));
SW0 switch1904 (.gate(net1083), .cc(\PD-xxxx10x0 ));
SW0 switch1905 (.gate(DBNeg), .cc(net648));
SW0 switch1906 (.gate(s7), .cc(net548));
SW0 switch1907 (.gate(net1020), .cc(net1277));
SW0 switch1908 (.gate(pipeUNK03), .cc(net1723));
SW0 switch1909 (.gate(pipeUNK03), .cc(net1614));
SW switch1910 (.gate(net1184), .cc1(net1631), .cc2(net903));
SW1 switch1911 (.gate(cclk), .cc(adh2));
SW switch1912 (.gate(net372), .cc1(net1085), .cc2(net1172));
SW switch1913 (.gate(notRdy0), .cc1(net912), .cc2(net1290));
SW0 switch1914 (.gate(\op-T2-abs-access ), .cc(net773));
SW0 switch1915 (.gate(net964), .cc(net17));
SW0 switch1916 (.gate(net964), .cc(clock1));
SW0 switch1917 (.gate(net663), .cc(\~pchp7 ));
SW0 switch1918 (.gate(net470), .cc(net1286));
SW0 switch1919 (.gate(net127), .cc(net135));
SW0 switch1920 (.gate(alu1), .cc(\~DA-ADD1 ));
SW switch1921 (.gate(net1245), .cc1(net299), .cc2(net1723));
SW1 switch1922 (.gate(net1152), .cc(ab2));
SW1 switch1923 (.gate(net1152), .cc(ab2));
SW1 switch1924 (.gate(net1152), .cc(ab2));
SW1 switch1925 (.gate(net1152), .cc(ab2));
SW1 switch1926 (.gate(net1152), .cc(ab2));
SW0 switch1927 (.gate(net1560), .cc(net1081));
SW0 switch1928 (.gate(net1609), .cc(ir5));
SW0 switch1929 (.gate(net1450), .cc(net1499));
SW0 switch1930 (.gate(RESG), .cc(net1712));
SW switch1931 (.gate(net1170), .cc1(net661), .cc2(net566));
SW switch1932 (.gate(cclk), .cc1(\~pclp5 ), .cc2(net1073));
SW0 switch1933 (.gate(net466), .cc(net7));
SW1 switch1934 (.gate(net466), .cc(net471));
SW0 switch1935 (.gate(net1258), .cc(net384));
SW0 switch1936 (.gate(\(AxB)2.~C12 ), .cc(\~(AxBxC)2 ));
SW0 switch1937 (.gate(\~ABH6 ), .cc(abh6));
SW switch1938 (.gate(cclk), .cc1(net1358), .cc2(net521));
SW0 switch1939 (.gate(net318), .cc(Pout1));
SW1 switch1940 (.gate(net1545), .cc(ab10));
SW switch1941 (.gate(cp1), .cc1(net644), .cc2(net428));
SW0 switch1942 (.gate(clk0), .cc(net519));
SW0 switch1943 (.gate(net1574), .cc(net1089));
SW0 switch1944 (.gate(\op-T5-jsr ), .cc(net1219));
SW0 switch1945 (.gate(y3), .cc(noty3));
SW0 switch1946 (.gate(net1411), .cc(\~pclp2 ));
SW0 switch1947 (.gate(net849), .cc(dpc33_PCHDB));
SW0 switch1948 (.gate(net862), .cc(net1211));
SW0 switch1949 (.gate(net94), .cc(net1024));
SW0 switch1950 (.gate(net933), .cc(net877));
SW switch1951 (.gate(net523), .cc1(net1657), .cc2(net1406));
SW switch1952 (.gate(net523), .cc1(net875), .cc2(net1659));
SW0 switch1953 (.gate(net523), .cc(net743));
SW0 switch1954 (.gate(\op-T+-bit ), .cc(net513));
SW0 switch1955 (.gate(net1230), .cc(net708));
SW1 switch1956 (.gate(net1230), .cc(dpc11_SBADD));
SW switch1957 (.gate(dpc13_ORS), .cc1(\~aluresult7 ), .cc2(\~(A+B)7 ));
SW switch1958 (.gate(dpc13_ORS), .cc1(\~(A+B)0 ), .cc2(\~aluresult0 ));
SW0 switch1959 (.gate(net947), .cc(net1654));
SW0 switch1960 (.gate(pcl6), .cc(net232));
SW switch1961 (.gate(dpc5_SADL), .cc1(adl0), .cc2(net332));
SW0 switch1962 (.gate(pd0), .cc(\pd0.clearIR ));
SW0 switch1963 (.gate(s2), .cc(net1190));
SW switch1964 (.gate(cclk), .cc1(net1300), .cc2(notir2));
SW switch1965 (.gate(net270), .cc1(net922), .cc2(BRtaken));
SW0 switch1966 (.gate(net270), .cc(net1115));
SW0 switch1967 (.gate(\~(A+B)2 ), .cc(\A+B2 ));
SW0 switch1968 (.gate(\~(A+B)2 ), .cc(C23));
SW0 switch1969 (.gate(\~pclp3 ), .cc(pclp3));
SW0 switch1970 (.gate(dor1), .cc(net794));
SW0 switch1971 (.gate(dor1), .cc(net288));
SW0 switch1972 (.gate(\op-shift ), .cc(net1681));
SW0 switch1973 (.gate(net43), .cc(net1270));
SW0 switch1974 (.gate(net1247), .cc(dpc39_PCLPCL));
SW0 switch1975 (.gate(net119), .cc(ir1));
SW switch1976 (.gate(C56), .cc1(net1390), .cc2(\~(AxBxC)6 ));
SW0 switch1977 (.gate(C56), .cc(\(AxB)6.~C56 ));
SW0 switch1978 (.gate(net188), .cc(t4));
SW switch1979 (.gate(net1303), .cc1(net782), .cc2(net1040));
SW0 switch1980 (.gate(adh4), .cc(net212));
SW0 switch1981 (.gate(pipephi2Reset0), .cc(net819));
SW0 switch1982 (.gate(idb3), .cc(net457));
SW0 switch1983 (.gate(net1033), .cc(dpc21_ADDADL));
SW switch1984 (.gate(dpc40_ADLPCL), .cc1(pcl7), .cc2(adl7));
SW switch1985 (.gate(dpc1_SBY), .cc1(y3), .cc2(sb3));
SW switch1986 (.gate(cclk), .cc1(net11), .cc2(net55));
SW0 switch1987 (.gate(net1274), .cc(net1069));
SW switch1988 (.gate(cp1), .cc1(net913), .cc2(net1274));
SW0 switch1989 (.gate(\op-T4-rti ), .cc(net604));
SW0 switch1990 (.gate(net23), .cc(net298));
SW1 switch1991 (.gate(net23), .cc(net1501));
SW0 switch1992 (.gate(net968), .cc(net1093));
SW switch1993 (.gate(cclk), .cc1(net1705), .cc2(net1020));
SW0 switch1994 (.gate(pipeUNK09), .cc(net781));
SW0 switch1995 (.gate(pipeUNK09), .cc(net1422));
SW0 switch1996 (.gate(net334), .cc(net118));
SW0 switch1997 (.gate(net700), .cc(net619));
SW0 switch1998 (.gate(\op-T2-stack-access ), .cc(net1090));
SW0 switch1999 (.gate(net1129), .cc(net1467));
SW1 switch2000 (.gate(net1633), .cc(ab5));
SW1 switch2001 (.gate(net1633), .cc(ab5));
SW1 switch2002 (.gate(net1633), .cc(ab5));
SW1 switch2003 (.gate(net1633), .cc(ab5));
SW1 switch2004 (.gate(net1633), .cc(ab5));
SW0 switch2005 (.gate(\~DA-ADD1 ), .cc(net1556));
SW0 switch2006 (.gate(\~DA-ADD1 ), .cc(net867));
SW0 switch2007 (.gate(net647), .cc(AxB5));
SW0 switch2008 (.gate(net1067), .cc(\ADH/ABH ));
SW switch2009 (.gate(cclk), .cc1(net541), .cc2(notir7));
SW switch2010 (.gate(cp1), .cc1(net1409), .cc2(net916));
SW0 switch2011 (.gate(net666), .cc(net862));
SW0 switch2012 (.gate(net1323), .cc(dpc37_PCLDB));
SW0 switch2013 (.gate(\~pchp7 ), .cc(pchp7));
SW0 switch2014 (.gate(\short-circuit-idx-add ), .cc(net1215));
SW0 switch2015 (.gate(net201), .cc(net1433));
SW0 switch2016 (.gate(idb7), .cc(DBNeg));
SW0 switch2017 (.gate(idb7), .cc(DBZ));
SW0 switch2018 (.gate(net636), .cc(nnT2BR));
SW1 switch2019 (.gate(net855), .cc(ab0));
SW1 switch2020 (.gate(net855), .cc(ab0));
SW1 switch2021 (.gate(net855), .cc(ab0));
SW1 switch2022 (.gate(net855), .cc(ab0));
SW1 switch2023 (.gate(net855), .cc(ab0));
SW0 switch2024 (.gate(notRdy0), .cc(net1343));
SW0 switch2025 (.gate(net646), .cc(net202));
SW0 switch2026 (.gate(cclk), .cc(net881));
SW switch2027 (.gate(net1056), .cc1(net1080), .cc2(net739));
SW1 switch2028 (.gate(cclk), .cc(adh7));
SW0 switch2029 (.gate(net878), .cc(net631));
SW0 switch2030 (.gate(net916), .cc(\short-circuit-idx-add ));
SW0 switch2031 (.gate(nnT2BR), .cc(net272));
SW switch2032 (.gate(cclk), .cc1(net80), .cc2(net1333));
SW0 switch2033 (.gate(\pd2.clearIR ), .cc(net571));
SW0 switch2034 (.gate(\pd2.clearIR ), .cc(\PD-xxx010x1 ));
SW0 switch2035 (.gate(\pd2.clearIR ), .cc(\PD-xxxx10x0 ));
SW0 switch2036 (.gate(\pd2.clearIR ), .cc(\PD-1xx000x0 ));
SW0 switch2037 (.gate(notidl4), .cc(idl4));
SW0 switch2038 (.gate(notidl4), .cc(idl4));
SW0 switch2039 (.gate(notidl4), .cc(idl4));
SW0 switch2040 (.gate(net196), .cc(dpc5_SADL));
SW0 switch2041 (.gate(\op-T0-jsr ), .cc(net1058));
SW switch2042 (.gate(cp1), .cc1(net1039), .cc2(net24));
SW0 switch2043 (.gate(\op-rti/rts ), .cc(net1649));
SW0 switch2044 (.gate(\op-rti/rts ), .cc(net1377));
SW switch2045 (.gate(cclk), .cc1(net1101), .cc2(net190));
SW0 switch2046 (.gate(\DC78.phi2 ), .cc(notalucout));
SW switch2047 (.gate(cclk), .cc1(net993), .cc2(net20));
SW0 switch2048 (.gate(\op-T5-rts ), .cc(net726));
SW0 switch2049 (.gate(net1455), .cc(net1412));
SW0 switch2050 (.gate(net1346), .cc(net1296));
SW1 switch2051 (.gate(net1346), .cc(net359));
SW0 switch2052 (.gate(\op-T+-shift-a ), .cc(net1455));
SW switch2053 (.gate(dpc19_ADDSB7), .cc1(alu7), .cc2(sb7));
SW0 switch2054 (.gate(net847), .cc(net104));
SW0 switch2055 (.gate(\op-T+-ora/and/eor/adc ), .cc(net1455));
SW0 switch2056 (.gate(net676), .cc(ab9));
SW0 switch2057 (.gate(net676), .cc(ab9));
SW0 switch2058 (.gate(net676), .cc(ab9));
SW0 switch2059 (.gate(net676), .cc(ab9));
SW0 switch2060 (.gate(net676), .cc(ab9));
SW0 switch2061 (.gate(net676), .cc(ab9));
SW0 switch2062 (.gate(net676), .cc(ab9));
SW0 switch2063 (.gate(net748), .cc(AxB7));
SW1 switch2064 (.gate(net1296), .cc(ab11));
SW0 switch2065 (.gate(net785), .cc(net267));
SW1 switch2066 (.gate(net1028), .cc(RnWstretched));
SW0 switch2067 (.gate(net1159), .cc(dasb2));
SW0 switch2068 (.gate(\pipe~VEC ), .cc(net1578));
SW0 switch2069 (.gate(net238), .cc(net1215));
SW0 switch2070 (.gate(net969), .cc(dpc0_YSB));
SW0 switch2071 (.gate(net232), .cc(net585));
SW0 switch2072 (.gate(net232), .cc(dpc34_PCLC));
SW0 switch2073 (.gate(net232), .cc(net1316));
SW switch2074 (.gate(cclk), .cc1(net1177), .cc2(net1069));
SW0 switch2075 (.gate(abh0), .cc(net1315));
SW0 switch2076 (.gate(abh0), .cc(net381));
SW switch2077 (.gate(cclk), .cc1(pipeUNK13), .cc2(net1045));
SW0 switch2078 (.gate(VEC1), .cc(\~VEC ));
SW switch2079 (.gate(cclk), .cc1(net728), .cc2(pipeVectorA0));
SW0 switch2080 (.gate(net781), .cc(net160));
SW0 switch2081 (.gate(VEC1), .cc(net912));
SW switch2082 (.gate(cclk), .cc1(pipeUNK30), .cc2(net385));
SW0 switch2084 (.gate(net646), .cc(net470));
SW switch2085 (.gate(cclk), .cc1(net1194), .cc2(pipeUNK04));
SW0 switch2086 (.gate(a4), .cc(net556));
SW0 switch2087 (.gate(\op-T2-php/pha ), .cc(net368));
SW0 switch2088 (.gate(\op-T2-php/pha ), .cc(\~WR ));
SW0 switch2089 (.gate(net1121), .cc(net291));
SW0 switch2090 (.gate(noty5), .cc(net733));
SW switch2091 (.gate(cclk), .cc1(\~ABL1 ), .cc2(net66));
SW1 switch2092 (.gate(abh4), .cc(net475));
SW0 switch2093 (.gate(abh4), .cc(net1677));
SW0 switch2094 (.gate(abh4), .cc(net999));
SW switch2095 (.gate(cclk), .cc1(\~aluresult0 ), .cc2(notalu0));
SW0 switch2096 (.gate(C01), .cc(\~C01 ));
SW switch2097 (.gate(C01), .cc1(net1510), .cc2(\~C12 ));
SW0 switch2098 (.gate(net1447), .cc(net1175));
SW0 switch2099 (.gate(\~C78 ), .cc(alurawcout));
SW0 switch2100 (.gate(net959), .cc(net1154));
SW0 switch2101 (.gate(net171), .cc(ab7));
SW0 switch2102 (.gate(net171), .cc(ab7));
SW0 switch2103 (.gate(net171), .cc(ab7));
SW0 switch2104 (.gate(net171), .cc(ab7));
SW switch2105 (.gate(net345), .cc1(dasb3), .cc2(net1686));
SW0 switch2106 (.gate(net345), .cc(net1097));
SW0 switch2107 (.gate(noty1), .cc(net767));
SW switch2108 (.gate(cp1), .cc1(net1387), .cc2(idl5));
SW0 switch2109 (.gate(net815), .cc(\0/ADL2 ));
SW0 switch2110 (.gate(\op-T0-cli/sei ), .cc(net1065));
SW0 switch2111 (.gate(pd5), .cc(\pd5.clearIR ));
SW0 switch2112 (.gate(x1), .cc(notx1));
SW0 switch2113 (.gate(net1505), .cc(net830));
SW0 switch2114 (.gate(net757), .cc(net1030));
SW switch2115 (.gate(cp1), .cc1(net1718), .cc2(net671));
SW0 switch2116 (.gate(net192), .cc(net1130));
SW0 switch2117 (.gate(net1024), .cc(net1069));
SW switch2118 (.gate(cclk), .cc1(net1231), .cc2(pipeUNK21));
SW0 switch2119 (.gate(\~ABH0 ), .cc(abh0));
SW0 switch2120 (.gate(clk0), .cc(net358));
SW0 switch2121 (.gate(net1222), .cc(net1090));
SW0 switch2122 (.gate(\op-T0-iny/dey ), .cc(net1717));
SW switch2123 (.gate(dpc3_SBX), .cc1(x0), .cc2(dasb0));
SW switch2124 (.gate(\~A.B6 ), .cc1(\~(AxB)6 ), .cc2(net482));
SW0 switch2126 (.gate(net1579), .cc(net221));
SW switch2127 (.gate(H1x1), .cc1(Pout4), .cc2(idb4));
SW0 switch2128 (.gate(db6), .cc(net374));
SW switch2129 (.gate(H1x1), .cc1(Pout3), .cc2(idb3));
SW switch2130 (.gate(H1x1), .cc1(Pout6), .cc2(idb6));
SW0 switch2131 (.gate(net507), .cc(net279));
SW switch2132 (.gate(net507), .cc1(net186), .cc2(net1082));
SW switch2133 (.gate(cp1), .cc1(net961), .cc2(notdor5));
SW0 switch2134 (.gate(net200), .cc(net1486));
SW switch2135 (.gate(net200), .cc1(net293), .cc2(net1367));
SW0 switch2136 (.gate(net200), .cc(net57));
SW0 switch2137 (.gate(RnWstretched), .cc(net1501));
SW0 switch2138 (.gate(RnWstretched), .cc(net1501));
SW switch2139 (.gate(cclk), .cc1(net952), .cc2(net1509));
SW0 switch2140 (.gate(notdor0), .cc(dor0));
SW0 switch2141 (.gate(aluvout), .cc(net1245));
SW0 switch2142 (.gate(pipeUNK04), .cc(net1644));
SW0 switch2143 (.gate(net108), .cc(dpc16_EORS));
SW0 switch2144 (.gate(net850), .cc(net1446));
SW0 switch2145 (.gate(net850), .cc(\short-circuit-branch-add ));
SW switch2146 (.gate(cclk), .cc1(net1169), .cc2(x0));
SW switch2147 (.gate(cclk), .cc1(net588), .cc2(notidl7));
SW1 switch2148 (.gate(cclk), .cc(adh5));
SW1 switch2149 (.gate(cclk), .cc(adl6));
SW0 switch2150 (.gate(RESP), .cc(net14));
SW0 switch2151 (.gate(NMIP), .cc(\~NMIP ));
SW0 switch2152 (.gate(net1534), .cc(net763));
SW1 switch2153 (.gate(net1534), .cc(dpc8_nDBADD));
SW0 switch2154 (.gate(net69), .cc(net1045));
SW switch2155 (.gate(net36), .cc1(dasb1), .cc2(net1322));
SW0 switch2156 (.gate(net36), .cc(net735));
SW1 switch2157 (.gate(net417), .cc(sync));
SW1 switch2158 (.gate(net417), .cc(sync));
SW1 switch2159 (.gate(net417), .cc(sync));
SW1 switch2160 (.gate(net417), .cc(sync));
SW1 switch2161 (.gate(net417), .cc(sync));
SW1 switch2162 (.gate(net417), .cc(sync));
SW1 switch2163 (.gate(net417), .cc(sync));
SW0 switch2164 (.gate(nnT2BR), .cc(net1211));
SW0 switch2165 (.gate(nnT2BR), .cc(net1211));
SW0 switch2166 (.gate(net1286), .cc(net1211));
SW0 switch2167 (.gate(t4), .cc(\op-T4-rts ));
SW0 switch2168 (.gate(t4), .cc(\op-T4-brk/jsr ));
SW0 switch2169 (.gate(t4), .cc(\op-T4-rti ));
SW0 switch2170 (.gate(t4), .cc(\op-T4-ind-y ));
SW0 switch2171 (.gate(t4), .cc(\op-T4-ind-x ));
SW0 switch2172 (.gate(t4), .cc(\op-T4-abs-idx ));
SW0 switch2173 (.gate(t4), .cc(\op-T4 ));
SW0 switch2174 (.gate(t4), .cc(\x-op-T4-ind-y ));
SW0 switch2175 (.gate(t4), .cc(\op-T4-brk ));
SW0 switch2176 (.gate(t4), .cc(\op-T4-jmp ));
SW0 switch2177 (.gate(t4), .cc(\x-op-T4-rti ));
SW0 switch2178 (.gate(t4), .cc(\op-T4-mem-abs-idx ));
SW1 switch2179 (.gate(net1399), .cc(cp1));
SW0 switch2180 (.gate(net398), .cc(net321));
SW0 switch2181 (.gate(net43), .cc(net692));
SW0 switch2182 (.gate(net1293), .cc(net620));
SW0 switch2183 (.gate(net936), .cc(\~C12 ));
SW0 switch2184 (.gate(p3), .cc(net1194));
SW0 switch2185 (.gate(\~A.B3 ), .cc(net988));
SW0 switch2186 (.gate(net743), .cc(net875));
SW switch2187 (.gate(net743), .cc1(net545), .cc2(net609));
SW0 switch2188 (.gate(net743), .cc(net1547));
SW0 switch2189 (.gate(notx2), .cc(net1694));
SW switch2190 (.gate(dpc27_SBADH), .cc1(adh7), .cc2(sb7));
SW switch2191 (.gate(dpc27_SBADH), .cc1(sb6), .cc2(adh6));
SW switch2192 (.gate(dpc1_SBY), .cc1(y0), .cc2(dasb0));
SW switch2193 (.gate(dpc27_SBADH), .cc1(adh0), .cc2(dasb0));
SW0 switch2194 (.gate(cp1), .cc(net38));
SW0 switch2195 (.gate(cp1), .cc(net1247));
SW0 switch2196 (.gate(net1252), .cc(net882));
SW switch2197 (.gate(dpc27_SBADH), .cc1(adh4), .cc2(dasb4));
SW switch2198 (.gate(dpc27_SBADH), .cc1(adh3), .cc2(sb3));
SW switch2199 (.gate(dpc27_SBADH), .cc1(adh2), .cc2(sb2));
SW switch2200 (.gate(net761), .cc1(net233), .cc2(net970));
SW0 switch2201 (.gate(net761), .cc(net762));
SW0 switch2202 (.gate(\dpc18_~DAA ), .cc(DC34));
SW0 switch2203 (.gate(\~op-branch-bit6 ), .cc(net1293));
SW0 switch2204 (.gate(y6), .cc(noty6));
SW0 switch2205 (.gate(dor0), .cc(net1072));
SW0 switch2206 (.gate(dor0), .cc(net769));
SW0 switch2207 (.gate(net755), .cc(net1170));
SW1 switch2208 (.gate(net834), .cc(net102));
SW0 switch2209 (.gate(net75), .cc(dpc20_ADDSB06));
SW0 switch2210 (.gate(C45), .cc(\~C45 ));
SW switch2211 (.gate(C45), .cc1(\~C56 ), .cc2(net165));
SW switch2212 (.gate(dpc15_ANDS), .cc1(\~A.B0 ), .cc2(\~aluresult0 ));
SW switch2213 (.gate(dpc15_ANDS), .cc1(\~A.B1 ), .cc2(\~aluresult1 ));
SW switch2214 (.gate(dpc15_ANDS), .cc1(\~A.B2 ), .cc2(\~aluresult2 ));
SW switch2215 (.gate(dpc15_ANDS), .cc1(\~A.B3 ), .cc2(\~aluresult3 ));
SW switch2216 (.gate(dpc15_ANDS), .cc1(\~A.B4 ), .cc2(\~aluresult4 ));
SW switch2217 (.gate(dpc15_ANDS), .cc1(\~aluresult5 ), .cc2(\~A.B5 ));
SW switch2218 (.gate(dpc15_ANDS), .cc1(\~A.B6 ), .cc2(\~aluresult6 ));
SW switch2219 (.gate(dpc15_ANDS), .cc1(\~aluresult7 ), .cc2(\~A.B7 ));
SW switch2220 (.gate(net233), .cc1(net1205), .cc2(net569));
SW1 switch2221 (.gate(cclk), .cc(adl1));
SW1 switch2222 (.gate(net1191), .cc(ab6));
SW1 switch2223 (.gate(net1191), .cc(ab6));
SW1 switch2224 (.gate(net1191), .cc(ab6));
SW1 switch2225 (.gate(net1191), .cc(ab6));
SW0 switch2226 (.gate(net1499), .cc(net709));
SW1 switch2227 (.gate(net1499), .cc(\dpc18_~DAA ));
SW0 switch2228 (.gate(net1549), .cc(net929));
SW0 switch2229 (.gate(cclk), .cc(dpc40_ADLPCL));
SW0 switch2230 (.gate(cclk), .cc(dpc39_PCLPCL));
SW0 switch2231 (.gate(net31), .cc(net132));
SW0 switch2232 (.gate(\A+B4 ), .cc(net1583));
SW0 switch2233 (.gate(\~A.B6 ), .cc(net112));
SW0 switch2234 (.gate(net756), .cc(\branch-forward.phi1 ));
SW switch2235 (.gate(dpc26_ACDB), .cc1(net146), .cc2(idb0));
SW switch2236 (.gate(dpc26_ACDB), .cc1(net929), .cc2(idb1));
SW switch2237 (.gate(dpc26_ACDB), .cc1(net1618), .cc2(idb2));
SW switch2238 (.gate(dpc26_ACDB), .cc1(net1654), .cc2(idb3));
SW switch2239 (.gate(dpc26_ACDB), .cc1(idb4), .cc2(net1344));
SW switch2240 (.gate(dpc26_ACDB), .cc1(net831), .cc2(idb5));
SW switch2241 (.gate(dpc26_ACDB), .cc1(net326), .cc2(idb6));
SW switch2242 (.gate(dpc26_ACDB), .cc1(net1592), .cc2(idb7));
SW0 switch2243 (.gate(pd4), .cc(\pd4.clearIR ));
SW switch2244 (.gate(net1345), .cc1(net1542), .cc2(net1685));
SW0 switch2245 (.gate(net1345), .cc(net1568));
SW0 switch2246 (.gate(net1649), .cc(net795));
SW switch2247 (.gate(cp1), .cc1(net1180), .cc2(net1533));
SW0 switch2248 (.gate(s0), .cc(net983));
SW0 switch2249 (.gate(\~DBZ ), .cc(net580));
SW1 switch2250 (.gate(abh2), .cc(net1545));
SW0 switch2251 (.gate(abh2), .cc(net1034));
SW0 switch2252 (.gate(abh2), .cc(net994));
SW0 switch2253 (.gate(\op-T2-mem-zp ), .cc(net347));
SW switch2254 (.gate(dpc27_SBADH), .cc1(sb1), .cc2(adh1));
SW0 switch2255 (.gate(dpc12_0ADD), .cc(alua2));
SW0 switch2256 (.gate(net610), .cc(net582));
SW switch2257 (.gate(dpc0_YSB), .cc1(net1251), .cc2(sb7));
SW0 switch2258 (.gate(pcl0), .cc(net937));
SW switch2259 (.gate(cclk), .cc1(net1500), .cc2(net526));
SW switch2260 (.gate(dpc0_YSB), .cc1(net658), .cc2(dasb4));
SW0 switch2261 (.gate(net47), .cc(net603));
SW switch2262 (.gate(dpc0_YSB), .cc1(net518), .cc2(sb6));
SW switch2263 (.gate(dpc0_YSB), .cc1(net733), .cc2(sb5));
SW0 switch2264 (.gate(pch5), .cc(net499));
SW0 switch2265 (.gate(\op-T3-jsr ), .cc(net824));
SW0 switch2266 (.gate(net862), .cc(net445));
SW0 switch2267 (.gate(pipeUNK36), .cc(\short-circuit-idx-add ));
SW switch2268 (.gate(cp1), .cc1(net738), .cc2(net1519));
SW0 switch2269 (.gate(\op-from-x ), .cc(net734));
SW1 switch2270 (.gate(cclk), .cc(idb5));
SW0 switch2271 (.gate(net50), .cc(net629));
SW switch2272 (.gate(cclk), .cc1(net440), .cc2(pipeUNK39));
SW0 switch2273 (.gate(\op-T3-branch ), .cc(net1716));
SW0 switch2274 (.gate(\op-T3-branch ), .cc(\~op-T3-branch ));
SW0 switch2275 (.gate(\op-T0-jmp ), .cc(net256));
SW0 switch2276 (.gate(\~pclp4 ), .cc(pclp4));
SW switch2278 (.gate(cclk), .cc1(net927), .cc2(notir4));
SW0 switch2279 (.gate(net628), .cc(net1335));
SW1 switch2280 (.gate(net628), .cc(dpc24_ACSB));
SW switch2281 (.gate(cclk), .cc1(net616), .cc2(net460));
SW0 switch2282 (.gate(notir6), .cc(\op-T0-cpy/iny ));
SW0 switch2283 (.gate(notir6), .cc(\op-T0-dex ));
SW0 switch2284 (.gate(notir6), .cc(\op-T0-cpx/inx ));
SW0 switch2285 (.gate(notir6), .cc(\op-T+-dex ));
SW0 switch2286 (.gate(notir6), .cc(\op-T+-inx ));
SW0 switch2287 (.gate(notir6), .cc(\op-T4-rts ));
SW0 switch2288 (.gate(notir6), .cc(\op-T5-rti ));
SW0 switch2289 (.gate(notir6), .cc(\op-ror ));
SW0 switch2290 (.gate(notir6), .cc(\op-T0-eor ));
SW0 switch2291 (.gate(notir6), .cc(\op-jmp ));
SW0 switch2292 (.gate(notir6), .cc(\op-T4-rti ));
SW0 switch2293 (.gate(notir6), .cc(\op-inc/nop ));
SW0 switch2294 (.gate(notir6), .cc(\op-rti/rts ));
SW0 switch2295 (.gate(notir6), .cc(\op-T0-cpx/cpy/inx/iny ));
SW0 switch2296 (.gate(notir6), .cc(\op-T0-cmp ));
SW0 switch2297 (.gate(notir6), .cc(\op-T0-sbc ));
SW0 switch2298 (.gate(notir6), .cc(\op-T0-adc/sbc ));
SW0 switch2299 (.gate(notir6), .cc(\op-T3-jmp ));
SW0 switch2300 (.gate(notir6), .cc(\op-T+-adc/sbc ));
SW0 switch2301 (.gate(notir6), .cc(\op-T0-pla ));
SW0 switch2302 (.gate(notir6), .cc(\op-T2-pha ));
SW0 switch2303 (.gate(notir6), .cc(\op-T0-shift-right-a ));
SW0 switch2304 (.gate(notir6), .cc(\op-shift-right ));
SW0 switch2305 (.gate(notir6), .cc(\op-T5-rts ));
SW0 switch2306 (.gate(notir6), .cc(\op-T0-jmp ));
SW0 switch2307 (.gate(notir6), .cc(\x-op-jmp ));
SW0 switch2308 (.gate(notir6), .cc(\op-T4-jmp ));
SW0 switch2309 (.gate(notir6), .cc(\op-T5-rti/rts ));
SW0 switch2310 (.gate(notir6), .cc(\op-T2-jmp-abs ));
SW0 switch2311 (.gate(notir6), .cc(\op-lsr/ror/dec/inc ));
SW0 switch2312 (.gate(notir6), .cc(\op-T0-cli/sei ));
SW0 switch2313 (.gate(notir6), .cc(\x-op-T+-adc/sbc ));
SW0 switch2314 (.gate(notir6), .cc(\x-op-T4-rti ));
SW0 switch2315 (.gate(notir6), .cc(\op-T+-cmp ));
SW0 switch2316 (.gate(notir6), .cc(\op-T+-cpx/cpy-abs ));
SW0 switch2317 (.gate(notir6), .cc(\op-T+-cpx/cpy-imm/zp ));
SW0 switch2318 (.gate(notir6), .cc(\op-T0-cld/sed ));
SW0 switch2319 (.gate(\~A.B2 ), .cc(net716));
SW switch2320 (.gate(dpc37_PCLDB), .cc1(pclp5), .cc2(idb5));
SW0 switch2321 (.gate(\~(A+B)0 ), .cc(\A+B0 ));
SW0 switch2322 (.gate(\~(A+B)0 ), .cc(C01));
SW0 switch2323 (.gate(\op-T3-stack/bit/jmp ), .cc(net604));
SW switch2324 (.gate(cclk), .cc1(net1455), .cc2(net1505));
SW0 switch2325 (.gate(net1566), .cc(net1240));
SW1 switch2326 (.gate(net1566), .cc(\dpc43_DL/DB ));
SW switch2327 (.gate(cp1), .cc1(net1507), .cc2(net864));
SW0 switch2328 (.gate(net1133), .cc(irline3));
SW switch2329 (.gate(dpc34_PCLC), .cc1(net856), .cc2(net919));
SW0 switch2330 (.gate(dpc34_PCLC), .cc(net835));
SW0 switch2331 (.gate(net581), .cc(net838));
SW switch2332 (.gate(net397), .cc1(net11), .cc2(net1563));
SW0 switch2333 (.gate(\op-brk/rti ), .cc(net134));
SW switch2334 (.gate(dpc37_PCLDB), .cc1(idb4), .cc2(pclp4));
SW0 switch2335 (.gate(net862), .cc(net1130));
SW1 switch2336 (.gate(cclk), .cc(adh3));
SW0 switch2337 (.gate(cclk), .cc(net133));
SW0 switch2338 (.gate(cclk), .cc(net161));
SW0 switch2339 (.gate(nots0), .cc(net332));
SW switch2340 (.gate(cclk), .cc1(\~aluresult2 ), .cc2(notalu2));
SW0 switch2341 (.gate(\op-rol/ror ), .cc(net1000));
SW0 switch2342 (.gate(net1257), .cc(net753));
SW0 switch2343 (.gate(net1257), .cc(net711));
SW0 switch2344 (.gate(net1257), .cc(net569));
SW0 switch2345 (.gate(net24), .cc(net440));
SW0 switch2346 (.gate(y0), .cc(noty0));
SW0 switch2347 (.gate(\op-T3-abs-idx ), .cc(net1107));
SW switch2348 (.gate(cclk), .cc1(net795), .cc2(net360));
SW switch2349 (.gate(net739), .cc1(dasb6), .cc2(net1554));
SW0 switch2350 (.gate(net739), .cc(net479));
SW switch2351 (.gate(cclk), .cc1(\~pclp3 ), .cc2(net1631));
SW0 switch2352 (.gate(\op-T5-rts ), .cc(net272));
SW1 switch2353 (.gate(net298), .cc(db7));
SW1 switch2354 (.gate(net298), .cc(db7));
SW1 switch2355 (.gate(net298), .cc(db7));
SW1 switch2356 (.gate(net298), .cc(db7));
SW0 switch2357 (.gate(net659), .cc(ab15));
SW0 switch2358 (.gate(net659), .cc(ab15));
SW0 switch2359 (.gate(net659), .cc(ab15));
SW0 switch2360 (.gate(net659), .cc(ab15));
SW0 switch2361 (.gate(net659), .cc(ab15));
SW0 switch2362 (.gate(net659), .cc(ab15));
SW switch2363 (.gate(dpc24_ACSB), .cc1(dasb0), .cc2(net146));
SW switch2364 (.gate(dpc24_ACSB), .cc1(sb1), .cc2(net929));
SW switch2365 (.gate(dpc24_ACSB), .cc1(net1618), .cc2(sb2));
SW switch2366 (.gate(dpc24_ACSB), .cc1(sb3), .cc2(net1654));
SW switch2367 (.gate(dpc24_ACSB), .cc1(dasb4), .cc2(net1344));
SW switch2368 (.gate(dpc24_ACSB), .cc1(sb5), .cc2(net831));
SW switch2369 (.gate(dpc24_ACSB), .cc1(net326), .cc2(sb6));
SW switch2370 (.gate(dpc24_ACSB), .cc1(net1592), .cc2(sb7));
SW switch2371 (.gate(dpc5_SADL), .cc1(adl1), .cc2(net694));
SW switch2372 (.gate(cclk), .cc1(\~ABL2 ), .cc2(net642));
SW0 switch2373 (.gate(\~pchp0 ), .cc(pchp0));
SW0 switch2374 (.gate(\dpc36_~IPC ), .cc(dpc34_PCLC));
SW0 switch2375 (.gate(notir3), .cc(\op-T2-abs-y ));
SW0 switch2376 (.gate(notir3), .cc(\op-T0-iny/dey ));
SW0 switch2377 (.gate(notir3), .cc(\x-op-T0-tya ));
SW0 switch2378 (.gate(notir3), .cc(\x-op-T0-txa ));
SW0 switch2379 (.gate(notir3), .cc(\op-T0-dex ));
SW0 switch2380 (.gate(notir3), .cc(\op-T0-txs ));
SW0 switch2381 (.gate(notir3), .cc(\op-T+-dex ));
SW0 switch2382 (.gate(notir3), .cc(\op-T+-inx ));
SW0 switch2383 (.gate(notir3), .cc(\op-T0-tsx ));
SW0 switch2384 (.gate(notir3), .cc(\op-T+-iny/dey ));
SW0 switch2385 (.gate(notir3), .cc(\op-T0-php/pha ));
SW0 switch2386 (.gate(notir3), .cc(\op-T3-plp/pla ));
SW0 switch2387 (.gate(notir3), .cc(\op-jmp ));
SW0 switch2388 (.gate(notir3), .cc(\op-T2-abs ));
SW0 switch2389 (.gate(notir3), .cc(\op-T3-abs-idx ));
SW0 switch2390 (.gate(notir3), .cc(\op-plp/pla ));
SW0 switch2391 (.gate(notir3), .cc(\op-T3-jmp ));
SW0 switch2392 (.gate(notir3), .cc(\op-T0-tya ));
SW0 switch2393 (.gate(notir3), .cc(\op-T+-shift-a ));
SW0 switch2394 (.gate(notir3), .cc(\op-T0-txa ));
SW0 switch2395 (.gate(notir3), .cc(\op-T0-pla ));
SW0 switch2396 (.gate(notir3), .cc(\op-T0-tay ));
SW0 switch2397 (.gate(notir3), .cc(\op-T0-shift-a ));
SW0 switch2398 (.gate(notir3), .cc(\op-T0-tax ));
SW0 switch2399 (.gate(notir3), .cc(\op-T4-abs-idx ));
SW0 switch2400 (.gate(notir3), .cc(\op-T2-pha ));
SW0 switch2401 (.gate(notir3), .cc(\op-T0-shift-right-a ));
SW0 switch2402 (.gate(notir3), .cc(\op-T2-abs-access ));
SW0 switch2403 (.gate(notir3), .cc(\op-T0-jmp ));
SW0 switch2404 (.gate(notir3), .cc(\op-T3-abs/idx/ind ));
SW0 switch2405 (.gate(notir3), .cc(\x-op-T3-abs-idx ));
SW0 switch2406 (.gate(notir3), .cc(\x-op-jmp ));
SW0 switch2407 (.gate(notir3), .cc(\op-push/pull ));
SW0 switch2408 (.gate(notir3), .cc(\op-T2-php ));
SW0 switch2409 (.gate(notir3), .cc(\op-T2-php/pha ));
SW0 switch2410 (.gate(notir3), .cc(\op-T4-jmp ));
SW0 switch2411 (.gate(notir3), .cc(\op-T2-jmp-abs ));
SW0 switch2412 (.gate(notir3), .cc(\x-op-T3-plp/pla ));
SW0 switch2413 (.gate(notir3), .cc(\op-T0-cli/sei ));
SW0 switch2414 (.gate(notir3), .cc(\op-T0-clc/sec ));
SW0 switch2415 (.gate(notir3), .cc(\op-T0-plp ));
SW0 switch2416 (.gate(notir3), .cc(\op-implied ));
SW0 switch2417 (.gate(notir3), .cc(\op-clv ));
SW0 switch2418 (.gate(notir3), .cc(\op-T+-cpx/cpy-abs ));
SW0 switch2419 (.gate(notir3), .cc(\op-T4-mem-abs-idx ));
SW0 switch2420 (.gate(notir3), .cc(\op-T+-asl/rol-a ));
SW0 switch2421 (.gate(notir3), .cc(\op-T3-mem-abs ));
SW0 switch2422 (.gate(notir3), .cc(\op-T0-cld/sed ));
SW0 switch2423 (.gate(notir3), .cc(\x-op-push/pull ));
SW0 switch2424 (.gate(net1255), .cc(dpc13_ORS));
SW0 switch2425 (.gate(net781), .cc(net1546));
SW0 switch2426 (.gate(net781), .cc(net1457));
SW0 switch2427 (.gate(net897), .cc(net1369));
SW0 switch2428 (.gate(net46), .cc(net1508));
SW0 switch2429 (.gate(alua5), .cc(net1559));
SW0 switch2430 (.gate(alua5), .cc(\~(A+B)5 ));
SW0 switch2431 (.gate(\op-rmw ), .cc(net510));
SW0 switch2432 (.gate(net1247), .cc(dpc40_ADLPCL));
SW0 switch2433 (.gate(net630), .cc(net152));
SW0 switch2434 (.gate(\~(AxB)2 ), .cc(net1572));
SW0 switch2435 (.gate(\~(AxB)2 ), .cc(\(AxB)2.~C12 ));
SW0 switch2436 (.gate(net335), .cc(\~WR ));
SW0 switch2437 (.gate(net1696), .cc(rw));
SW0 switch2438 (.gate(net1696), .cc(rw));
SW0 switch2439 (.gate(net1696), .cc(rw));
SW0 switch2440 (.gate(net1696), .cc(rw));
SW0 switch2441 (.gate(net1696), .cc(rw));
SW0 switch2442 (.gate(dpc28_0ADH0), .cc(adh0));
SW0 switch2443 (.gate(net192), .cc(net506));
SW0 switch2444 (.gate(\op-store ), .cc(\~op-store ));
SW0 switch2445 (.gate(\op-SRS ), .cc(net139));
SW switch2446 (.gate(cclk), .cc1(nots1), .cc2(net1711));
SW1 switch2447 (.gate(net1545), .cc(ab10));
SW switch2448 (.gate(net754), .cc1(net648), .cc2(net1181));
SW0 switch2449 (.gate(net754), .cc(net1595));
SW switch2450 (.gate(dpc30_ADHPCH), .cc1(pch1), .cc2(adh1));
SW switch2451 (.gate(cp1), .cc1(net590), .cc2(net1178));
SW0 switch2452 (.gate(\~ABH5 ), .cc(abh5));
SW switch2453 (.gate(dpc30_ADHPCH), .cc1(pch0), .cc2(adh0));
SW0 switch2454 (.gate(abh1), .cc(net617));
SW0 switch2455 (.gate(abh1), .cc(net676));
SW switch2456 (.gate(cclk), .cc1(\~pchp6 ), .cc2(net1192));
SW1 switch2457 (.gate(abh7), .cc(net1639));
SW0 switch2458 (.gate(abh7), .cc(net1153));
SW0 switch2459 (.gate(abh7), .cc(net659));
SW0 switch2460 (.gate(net1018), .cc(net100));
SW0 switch2461 (.gate(AxB5), .cc(\~(AxB)5 ));
SW0 switch2462 (.gate(net231), .cc(ONEBYTE));
SW0 switch2463 (.gate(\x-op-T3-plp/pla ), .cc(net368));
SW0 switch2464 (.gate(net877), .cc(net911));
SW0 switch2465 (.gate(net877), .cc(net911));
SW0 switch2466 (.gate(net300), .cc(net847));
SW0 switch2467 (.gate(net133), .cc(net602));
SW1 switch2468 (.gate(net133), .cc(dpc2_XSB));
SW0 switch2469 (.gate(net709), .cc(\dpc18_~DAA ));
SW0 switch2470 (.gate(x0), .cc(notx0));
SW0 switch2471 (.gate(net318), .cc(net1293));
SW0 switch2472 (.gate(db4), .cc(net1075));
SW0 switch2473 (.gate(dpc34_PCLC), .cc(net1007));
SW0 switch2474 (.gate(net236), .cc(net176));
SW switch2475 (.gate(dpc31_PCHPCH), .cc1(pch6), .cc2(pchp6));
SW switch2476 (.gate(dpc31_PCHPCH), .cc1(pch7), .cc2(pchp7));
SW switch2477 (.gate(dpc31_PCHPCH), .cc1(pch4), .cc2(pchp4));
SW switch2478 (.gate(dpc31_PCHPCH), .cc1(pch5), .cc2(pchp5));
SW switch2479 (.gate(dpc31_PCHPCH), .cc1(pch2), .cc2(pchp2));
SW switch2480 (.gate(dpc31_PCHPCH), .cc1(pch3), .cc2(pchp3));
SW switch2481 (.gate(dpc31_PCHPCH), .cc1(pch0), .cc2(pchp0));
SW switch2482 (.gate(dpc31_PCHPCH), .cc1(pch1), .cc2(pchp1));
SW switch2483 (.gate(cclk), .cc1(net515), .cc2(net1411));
SW0 switch2484 (.gate(\op-T0-ldy-mem ), .cc(net616));
SW0 switch2485 (.gate(dpc29_0ADH17), .cc(adh3));
SW0 switch2486 (.gate(dpc29_0ADH17), .cc(adh2));
SW0 switch2487 (.gate(dpc29_0ADH17), .cc(adh5));
SW0 switch2488 (.gate(dpc29_0ADH17), .cc(adh4));
SW0 switch2489 (.gate(\op-ANDS ), .cc(net550));
SW0 switch2490 (.gate(dpc29_0ADH17), .cc(adh7));
SW0 switch2491 (.gate(dpc29_0ADH17), .cc(adh6));
SW0 switch2492 (.gate(net360), .cc(net1230));
SW0 switch2493 (.gate(\op-T2-ADL/ADD ), .cc(net1118));
SW switch2494 (.gate(net1289), .cc1(net632), .cc2(net1058));
SW0 switch2495 (.gate(pipeUNK37), .cc(net198));
SW0 switch2496 (.gate(pipeUNK37), .cc(net198));
SW0 switch2497 (.gate(\~IRQP ), .cc(net1092));
SW switch2498 (.gate(fetch), .cc1(net1675), .cc2(net74));
SW switch2499 (.gate(fetch), .cc1(net1609), .cc2(net1378));
SW switch2500 (.gate(net270), .cc1(net1692), .cc2(net1082));
SW0 switch2501 (.gate(adh0), .cc(net1668));
SW0 switch2502 (.gate(\op-T2-brk ), .cc(net824));
SW switch2503 (.gate(dpc8_nDBADD), .cc1(alub1), .cc2(net583));
SW switch2504 (.gate(dpc8_nDBADD), .cc1(alub3), .cc2(net1621));
SW0 switch2505 (.gate(net182), .cc(net1619));
SW switch2506 (.gate(cclk), .cc1(net126), .cc2(net1486));
SW0 switch2507 (.gate(\op-T2 ), .cc(net152));
SW0 switch2508 (.gate(pipeUNK02), .cc(net1492));
SW0 switch2509 (.gate(net1357), .cc(net378));
SW0 switch2510 (.gate(net1161), .cc(net732));
SW0 switch2511 (.gate(idb3), .cc(net1621));
SW0 switch2512 (.gate(net646), .cc(net182));
SW0 switch2513 (.gate(\op-T3-mem-abs ), .cc(net347));
SW switch2514 (.gate(cp1), .cc1(net1267), .cc2(net1298));
SW0 switch2515 (.gate(net1613), .cc(net42));
SW1 switch2516 (.gate(net1613), .cc(net643));
SW0 switch2517 (.gate(\~DA-ADD1 ), .cc(net1682));
SW0 switch2518 (.gate(\~DA-ADD1 ), .cc(net1362));
SW switch2519 (.gate(cclk), .cc1(pipeT5out), .cc2(net378));
SW0 switch2520 (.gate(notRdy0), .cc(notRnWprepad));
SW0 switch2521 (.gate(notRdy0), .cc(net1718));
SW0 switch2522 (.gate(\op-T0-eor ), .cc(net837));
SW1 switch2523 (.gate(net747), .cc(clk1out));
SW0 switch2524 (.gate(net358), .cc(net1715));
SW switch2525 (.gate(dpc38_PCLADL), .cc1(adl4), .cc2(pclp4));
SW switch2526 (.gate(dpc38_PCLADL), .cc1(pclp5), .cc2(adl5));
SW switch2527 (.gate(dpc38_PCLADL), .cc1(adl6), .cc2(pclp6));
SW switch2528 (.gate(dpc38_PCLADL), .cc1(pclp7), .cc2(adl7));
SW switch2529 (.gate(dpc38_PCLADL), .cc1(adl0), .cc2(pclp0));
SW switch2530 (.gate(dpc38_PCLADL), .cc1(pclp1), .cc2(adl1));
SW switch2531 (.gate(dpc38_PCLADL), .cc1(adl2), .cc2(pclp2));
SW switch2532 (.gate(dpc38_PCLADL), .cc1(pclp3), .cc2(adl3));
SW0 switch2533 (.gate(net854), .cc(net975));
SW0 switch2534 (.gate(net1345), .cc(net1500));
SW switch2535 (.gate(cclk), .cc1(net635), .cc2(\~ABH6 ));
SW0 switch2536 (.gate(net1404), .cc(net133));
SW0 switch2537 (.gate(\0/ADL2 ), .cc(adl2));
SW0 switch2538 (.gate(idb6), .cc(net1416));
SW0 switch2539 (.gate(net1276), .cc(net930));
SW0 switch2540 (.gate(net1276), .cc(net930));
SW0 switch2541 (.gate(net1400), .cc(net83));
SW0 switch2542 (.gate(net1509), .cc(net611));
SW0 switch2543 (.gate(adl3), .cc(net1507));
SW1 switch2544 (.gate(net839), .cc(net43));
SW switch2545 (.gate(cclk), .cc1(net484), .cc2(\~pclp7 ));
SW0 switch2546 (.gate(net43), .cc(net6));
SW switch2547 (.gate(dpc32_PCHADH), .cc1(adh7), .cc2(pchp7));
SW switch2548 (.gate(dpc32_PCHADH), .cc1(adh6), .cc2(pchp6));
SW switch2549 (.gate(dpc32_PCHADH), .cc1(adh5), .cc2(pchp5));
SW switch2550 (.gate(dpc32_PCHADH), .cc1(adh4), .cc2(pchp4));
SW switch2551 (.gate(dpc32_PCHADH), .cc1(adh3), .cc2(pchp3));
SW switch2552 (.gate(dpc32_PCHADH), .cc1(adh2), .cc2(pchp2));
SW switch2553 (.gate(dpc32_PCHADH), .cc1(adh1), .cc2(pchp1));
SW switch2554 (.gate(dpc32_PCHADH), .cc1(adh0), .cc2(pchp0));
SW switch2555 (.gate(net1440), .cc1(net605), .cc2(net779));
SW0 switch2556 (.gate(\dpc18_~DAA ), .cc(net700));
SW switch2557 (.gate(cclk), .cc1(\~ABH0 ), .cc2(net381));
SW0 switch2558 (.gate(cp1), .cc(net1129));
SW0 switch2559 (.gate(net1642), .cc(\~WR ));
SW1 switch2560 (.gate(net1041), .cc(ab3));
SW1 switch2561 (.gate(net1041), .cc(ab3));
SW1 switch2562 (.gate(net1041), .cc(ab3));
SW1 switch2563 (.gate(net1041), .cc(ab3));
SW1 switch2564 (.gate(net1041), .cc(ab3));
SW0 switch2565 (.gate(abl6), .cc(net1254));
SW0 switch2566 (.gate(abl6), .cc(net1195));
SW1 switch2567 (.gate(abl6), .cc(net1191));
SW0 switch2568 (.gate(net389), .cc(net300));
SW0 switch2569 (.gate(net1541), .cc(net491));
SW1 switch2570 (.gate(net1541), .cc(dpc10_ADLADD));
SW0 switch2571 (.gate(cclk), .cc(net431));
SW1 switch2572 (.gate(net1639), .cc(ab15));
SW1 switch2573 (.gate(net475), .cc(ab12));
SW0 switch2574 (.gate(RnWstretched), .cc(net1072));
SW0 switch2575 (.gate(RnWstretched), .cc(net1072));
SW0 switch2576 (.gate(pipeUNK29), .cc(net1189));
SW0 switch2577 (.gate(pipeUNK29), .cc(net1511));
SW switch2578 (.gate(net410), .cc1(net344), .cc2(net814));
SW0 switch2579 (.gate(net410), .cc(net557));
SW0 switch2580 (.gate(\~(AxB)4 ), .cc(net375));
SW0 switch2581 (.gate(\~(AxB)4 ), .cc(\(AxB)4.~C34 ));
SW switch2582 (.gate(cclk), .cc1(pipeT3out), .cc2(net678));
SW0 switch2583 (.gate(pipeUNK22), .cc(net533));
SW0 switch2584 (.gate(net410), .cc(net474));
SW0 switch2585 (.gate(net1423), .cc(net1608));
SW1 switch2586 (.gate(net1423), .cc(net869));
SW switch2587 (.gate(cp1), .cc1(net168), .cc2(net836));
SW0 switch2588 (.gate(nmi), .cc(net1392));
SW switch2589 (.gate(cclk), .cc1(net1699), .cc2(net1024));
SW0 switch2590 (.gate(\~ABL4 ), .cc(abl4));
SW switch2591 (.gate(cp1), .cc1(net468), .cc2(net18));
SW switch2592 (.gate(dpc13_ORS), .cc1(\~(A+B)4 ), .cc2(\~aluresult4 ));
SW0 switch2593 (.gate(net389), .cc(net1649));
SW0 switch2594 (.gate(\op-T3-plp/pla ), .cc(net1464));
SW switch2595 (.gate(dpc13_ORS), .cc1(\~(A+B)5 ), .cc2(\~aluresult5 ));
SW0 switch2596 (.gate(net18), .cc(net378));
SW switch2597 (.gate(net1570), .cc1(net1480), .cc2(\dpc36_~IPC ));
SW1 switch2598 (.gate(cclk), .cc(idb6));
SW switch2599 (.gate(net440), .cc1(net1681), .cc2(net905));
SW switch2600 (.gate(cclk), .cc1(net213), .cc2(notidl1));
SW switch2601 (.gate(cclk), .cc1(net862), .cc2(\pipeT-SYNC ));
SW switch2602 (.gate(cp1), .cc1(net789), .cc2(notdor7));
SW0 switch2603 (.gate(net1166), .cc(net1685));
SW0 switch2604 (.gate(net1166), .cc(net1568));
SW0 switch2605 (.gate(net1660), .cc(net855));
SW1 switch2606 (.gate(net1660), .cc(net1100));
SW0 switch2607 (.gate(\~VEC ), .cc(net1712));
SW0 switch2608 (.gate(\x-op-push/pull ), .cc(\op-implied ));
SW switch2609 (.gate(net779), .cc1(net656), .cc2(net1594));
SW0 switch2610 (.gate(\~NMIP ), .cc(NMIP));
SW0 switch2611 (.gate(net556), .cc(net1344));
SW0 switch2612 (.gate(\op-EORS ), .cc(\op-SUMS ));
SW0 switch2613 (.gate(net1315), .cc(net826));
SW0 switch2614 (.gate(net1265), .cc(net1202));
SW0 switch2615 (.gate(net1265), .cc(dpc35_PCHC));
SW switch2616 (.gate(cclk), .cc1(net733), .cc2(y5));
SW1 switch2617 (.gate(net1639), .cc(ab15));
SW0 switch2618 (.gate(notdor7), .cc(dor7));
SW0 switch2619 (.gate(pipeT4out), .cc(net1703));
SW0 switch2620 (.gate(pipeT4out), .cc(net395));
SW0 switch2621 (.gate(net1153), .cc(net1639));
SW1 switch2622 (.gate(net1153), .cc(net659));
SW0 switch2623 (.gate(alu5), .cc(net761));
SW0 switch2624 (.gate(net781), .cc(net1550));
SW switch2625 (.gate(cclk), .cc1(nnT2BR), .cc2(net1269));
SW0 switch2626 (.gate(\~(AxB)6 ), .cc(net1390));
SW0 switch2627 (.gate(\~(AxB)6 ), .cc(\(AxB)6.~C56 ));
SW0 switch2628 (.gate(\op-T0-shift-a ), .cc(net11));
SW switch2629 (.gate(cclk), .cc1(pipeUNK09), .cc2(net327));
SW switch2630 (.gate(cclk), .cc1(\~op-set-C ), .cc2(pipeUNK08));
SW switch2631 (.gate(cp1), .cc1(notRnWprepad), .cc2(net1579));
SW switch2632 (.gate(cp1), .cc1(p1), .cc2(net566));
SW0 switch2633 (.gate(net1247), .cc(dpc3_SBX));
SW switch2634 (.gate(cclk), .cc1(net306), .cc2(net581));
SW0 switch2635 (.gate(net1157), .cc(\dpc41_DL/ADL ));
SW0 switch2636 (.gate(net562), .cc(NMIL));
SW0 switch2637 (.gate(notdor5), .cc(dor5));
SW1 switch2638 (.gate(net1639), .cc(ab15));
SW0 switch2639 (.gate(idb2), .cc(DBZ));
SW0 switch2640 (.gate(notalu5), .cc(alu5));
SW0 switch2641 (.gate(idb2), .cc(net1573));
SW0 switch2642 (.gate(net625), .cc(net662));
SW1 switch2643 (.gate(net625), .cc(dpc3_SBX));
SW0 switch2644 (.gate(net646), .cc(net1172));
SW0 switch2645 (.gate(notidl3), .cc(idl3));
SW0 switch2646 (.gate(notidl3), .cc(idl3));
SW0 switch2647 (.gate(notidl3), .cc(idl3));
SW0 switch2648 (.gate(\~C12 ), .cc(C12));
SW0 switch2649 (.gate(\~C12 ), .cc(net433));
SW0 switch2650 (.gate(net609), .cc(net1213));
SW1 switch2651 (.gate(dor0), .cc(net1325));
SW0 switch2652 (.gate(net604), .cc(net385));
SW0 switch2653 (.gate(net1145), .cc(\op-ORS ));
SW0 switch2654 (.gate(a0), .cc(net5));
SW0 switch2655 (.gate(\op-T2-abs-y ), .cc(net1717));
SW switch2656 (.gate(cclk), .cc1(\pipe~T0 ), .cc2(net17));
SW0 switch2657 (.gate(pipeT5out), .cc(net1615));
SW0 switch2658 (.gate(net359), .cc(ab11));
SW0 switch2659 (.gate(net359), .cc(ab11));
SW0 switch2660 (.gate(net359), .cc(ab11));
SW0 switch2661 (.gate(net359), .cc(ab11));
SW0 switch2662 (.gate(net359), .cc(ab11));
SW0 switch2663 (.gate(net359), .cc(ab11));
SW0 switch2664 (.gate(net359), .cc(ab11));
SW0 switch2665 (.gate(net790), .cc(net191));
SW0 switch2666 (.gate(\op-T2-ind-y ), .cc(net1107));
SW0 switch2667 (.gate(db6), .cc(net1638));
SW switch2668 (.gate(\ADH/ABH ), .cc1(\~ABH2 ), .cc2(net836));
SW0 switch2669 (.gate(\~alucout ), .cc(\~~alucout ));
SW0 switch2670 (.gate(\xx-op-T5-jsr ), .cc(net368));
SW0 switch2671 (.gate(alua0), .cc(net316));
SW0 switch2672 (.gate(alua0), .cc(\~(A+B)0 ));
SW0 switch2673 (.gate(\0/ADL0 ), .cc(net696));
SW0 switch2674 (.gate(abl5), .cc(net210));
SW0 switch2675 (.gate(abl5), .cc(net172));
SW1 switch2676 (.gate(abl5), .cc(net1633));
SW0 switch2677 (.gate(net419), .cc(net1618));
SW0 switch2678 (.gate(cp1), .cc(net43));
SW0 switch2679 (.gate(cp1), .cc(net1247));
SW0 switch2680 (.gate(cp1), .cc(net1247));
SW0 switch2681 (.gate(a3), .cc(net947));
SW0 switch2682 (.gate(idb1), .cc(net243));
SW switch2683 (.gate(dpc9_DBADD), .cc1(alub7), .cc2(idb7));
SW switch2684 (.gate(dpc9_DBADD), .cc1(alub6), .cc2(idb6));
SW0 switch2685 (.gate(ir3), .cc(\op-T3-ind-y ));
SW0 switch2686 (.gate(ir3), .cc(\op-T2-ind-x ));
SW0 switch2687 (.gate(ir3), .cc(\op-T0-jsr ));
SW0 switch2688 (.gate(ir3), .cc(\op-T5-brk ));
SW0 switch2689 (.gate(ir3), .cc(\op-T4-rts ));
SW0 switch2690 (.gate(ir3), .cc(\op-T5-rti ));
SW0 switch2691 (.gate(ir3), .cc(\op-T2-ADL/ADD ));
SW0 switch2692 (.gate(ir3), .cc(\op-T4-brk/jsr ));
SW0 switch2693 (.gate(ir3), .cc(\op-T4-rti ));
SW0 switch2694 (.gate(ir3), .cc(\op-T3-ind-x ));
SW0 switch2695 (.gate(ir3), .cc(\op-T4-ind-y ));
SW0 switch2696 (.gate(ir3), .cc(\op-T2-ind-y ));
SW0 switch2697 (.gate(ir3), .cc(\op-T4-ind-x ));
SW0 switch2698 (.gate(ir3), .cc(\x-op-T3-ind-y ));
SW0 switch2699 (.gate(ir3), .cc(\op-rti/rts ));
SW0 switch2700 (.gate(ir3), .cc(\op-T2-jsr ));
SW0 switch2701 (.gate(ir3), .cc(\op-T5-jsr ));
SW0 switch2702 (.gate(ir3), .cc(\op-T5-ind-y ));
SW0 switch2703 (.gate(ir3), .cc(\op-branch-done ));
SW0 switch2704 (.gate(ir3), .cc(\op-T2-brk ));
SW0 switch2705 (.gate(ir3), .cc(\op-T3-jsr ));
SW0 switch2706 (.gate(ir3), .cc(\op-T2-branch ));
SW0 switch2707 (.gate(ir3), .cc(\op-T2-zp/zp-idx ));
SW0 switch2708 (.gate(ir3), .cc(\op-T2-ind ));
SW0 switch2709 (.gate(ir3), .cc(\op-T5-rts ));
SW0 switch2710 (.gate(ir3), .cc(\op-T0-brk/rti ));
SW0 switch2711 (.gate(ir3), .cc(\op-T5-ind-x ));
SW0 switch2712 (.gate(ir3), .cc(\x-op-T4-ind-y ));
SW0 switch2713 (.gate(ir3), .cc(\op-T3-branch ));
SW0 switch2714 (.gate(ir3), .cc(\op-brk/rti ));
SW0 switch2715 (.gate(ir3), .cc(\op-jsr ));
SW0 switch2716 (.gate(ir3), .cc(\op-T4-brk ));
SW0 switch2717 (.gate(ir3), .cc(\op-T5-rti/rts ));
SW0 switch2718 (.gate(ir3), .cc(\xx-op-T5-jsr ));
SW0 switch2719 (.gate(ir3), .cc(\op-T3-mem-zp-idx ));
SW0 switch2720 (.gate(ir3), .cc(\x-op-T4-rti ));
SW0 switch2721 (.gate(ir3), .cc(\op-T+-cpx/cpy-imm/zp ));
SW0 switch2722 (.gate(ir3), .cc(\op-T2-mem-zp ));
SW0 switch2723 (.gate(ir3), .cc(\op-T5-mem-ind-idx ));
SW switch2724 (.gate(cp1), .cc1(net1147), .cc2(idl7));
SW switch2725 (.gate(dpc9_DBADD), .cc1(alub1), .cc2(idb1));
SW switch2726 (.gate(dpc9_DBADD), .cc1(alub3), .cc2(idb3));
SW switch2727 (.gate(dpc9_DBADD), .cc1(idb2), .cc2(alub2));
SW switch2728 (.gate(dpc9_DBADD), .cc1(alub5), .cc2(idb5));
SW switch2729 (.gate(dpc9_DBADD), .cc1(alub4), .cc2(idb4));
SW switch2731 (.gate(cclk), .cc1(x5), .cc2(net578));
SW0 switch2732 (.gate(\op-T0-tsx ), .cc(net1586));
SW switch2733 (.gate(cclk), .cc1(\~ABH2 ), .cc2(net994));
SW switch2734 (.gate(net1316), .cc1(net1386), .cc2(net426));
SW0 switch2735 (.gate(net1316), .cc(net914));
SW1 switch2736 (.gate(cclk), .cc(adl0));
SW switch2737 (.gate(cclk), .cc1(net1229), .cc2(\~pchp0 ));
SW0 switch2738 (.gate(net1441), .cc(\dpc42_DL/ADH ));
SW switch2739 (.gate(alub7), .cc1(\~A.B7 ), .cc2(net1695));
SW0 switch2740 (.gate(alub7), .cc(\~(A+B)7 ));
SW0 switch2741 (.gate(net1316), .cc(net20));
SW0 switch2742 (.gate(net853), .cc(net387));
SW0 switch2743 (.gate(net519), .cc(net670));
SW0 switch2744 (.gate(net519), .cc(net670));
SW switch2745 (.gate(dpc37_PCLDB), .cc1(pclp3), .cc2(idb3));
SW switch2746 (.gate(dpc37_PCLDB), .cc1(pclp1), .cc2(idb1));
SW switch2747 (.gate(dpc37_PCLDB), .cc1(idb7), .cc2(pclp7));
SW0 switch2748 (.gate(net698), .cc(VEC1));
SW0 switch2749 (.gate(net846), .cc(net1371));
SW0 switch2750 (.gate(\dpc18_~DAA ), .cc(DC78));
SW0 switch2751 (.gate(net21), .cc(net228));
SW1 switch2752 (.gate(net21), .cc(dpc30_ADHPCH));
SW switch2753 (.gate(cclk), .cc1(pipeUNK01), .cc2(\branch-forward.phi1 ));
SW0 switch2754 (.gate(notalu7), .cc(alu7));
SW0 switch2755 (.gate(pipeUNK14), .cc(net661));
SW0 switch2756 (.gate(pipeUNK30), .cc(net1178));
SW switch2757 (.gate(cclk), .cc1(net1121), .cc2(net1225));
SW0 switch2758 (.gate(net1247), .cc(dpc11_SBADD));
SW0 switch2759 (.gate(pcl2), .cc(net783));
SW0 switch2760 (.gate(\pd4.clearIR ), .cc(net227));
SW0 switch2761 (.gate(net602), .cc(dpc2_XSB));
SW switch2762 (.gate(cp1), .cc1(net1661), .cc2(idl3));
SW0 switch2763 (.gate(net611), .cc(net255));
SW1 switch2764 (.gate(net611), .cc(dpc31_PCHPCH));
SW0 switch2765 (.gate(notRdy0), .cc(net917));
SW0 switch2766 (.gate(net954), .cc(net513));
SW0 switch2767 (.gate(net1026), .cc(net322));
SW1 switch2768 (.gate(net1026), .cc(net171));
SW switch2769 (.gate(pipeUNK16), .cc1(net455), .cc2(net1082));
SW switch2770 (.gate(DBNeg), .cc1(\branch-back ), .cc2(net1249));
SW switch2771 (.gate(cclk), .cc1(pipeUNK40), .cc2(net191));
SW0 switch2772 (.gate(\op-T+-adc/sbc ), .cc(net1455));
SW0 switch2773 (.gate(\~(A+B)4 ), .cc(\A+B4 ));
SW0 switch2774 (.gate(\~(A+B)4 ), .cc(C45));
SW0 switch2775 (.gate(cclk), .cc(dpc26_ACDB));
SW0 switch2776 (.gate(cclk), .cc(dpc24_ACSB));
SW0 switch2777 (.gate(net842), .cc(net1479));
SW1 switch2778 (.gate(net842), .cc(net66));
SW1 switch2779 (.gate(abh1), .cc(net1140));
SW0 switch2780 (.gate(net1409), .cc(net1231));
SW0 switch2781 (.gate(\op-ANDS ), .cc(net11));
SW0 switch2782 (.gate(sb5), .cc(net1135));
SW0 switch2783 (.gate(alua7), .cc(net1695));
SW0 switch2784 (.gate(alua7), .cc(\~(A+B)7 ));
SW switch2785 (.gate(cclk), .cc1(\~ABL4 ), .cc2(net86));
SW0 switch2786 (.gate(net70), .cc(net1117));
SW0 switch2787 (.gate(net1211), .cc(net10));
SW0 switch2788 (.gate(net637), .cc(notaluvout));
SW1 switch2789 (.gate(net1608), .cc(ab13));
SW switch2790 (.gate(net1599), .cc1(net807), .cc2(net431));
SW0 switch2791 (.gate(net1335), .cc(dpc24_ACSB));
SW0 switch2792 (.gate(\op-T+-asl/rol-a ), .cc(\~op-set-C ));
SW0 switch2793 (.gate(net1247), .cc(dpc2_XSB));
SW switch2794 (.gate(C67), .cc1(notaluvout), .cc2(net1489));
SW0 switch2795 (.gate(C67), .cc(net637));
SW0 switch2796 (.gate(pipeUNK23), .cc(net819));
SW0 switch2797 (.gate(noty4), .cc(net658));
SW switch2798 (.gate(dpc8_nDBADD), .cc1(alub5), .cc2(net1383));
SW switch2799 (.gate(dpc8_nDBADD), .cc1(alub6), .cc2(net351));
SW switch2800 (.gate(dpc8_nDBADD), .cc1(alub7), .cc2(net423));
SW0 switch2801 (.gate(net1605), .cc(\PD-1xx000x0 ));
SW0 switch2802 (.gate(net927), .cc(ir4));
SW0 switch2803 (.gate(net958), .cc(net1449));
SW switch2804 (.gate(cclk), .cc1(net871), .cc2(x7));
SW switch2805 (.gate(net919), .cc1(net1229), .cc2(net835));
SW switch2806 (.gate(net919), .cc1(net1486), .cc2(net1538));
SW0 switch2807 (.gate(net919), .cc(net200));
SW0 switch2808 (.gate(net1211), .cc(net1655));
SW0 switch2809 (.gate(clearIR), .cc(\pd1.clearIR ));
SW0 switch2810 (.gate(clearIR), .cc(\pd7.clearIR ));
SW switch2811 (.gate(cp1), .cc1(net705), .cc2(net1668));
SW0 switch2812 (.gate(\op-T2-abs-access ), .cc(net1211));
SW0 switch2813 (.gate(net1492), .cc(net1445));
SW0 switch2814 (.gate(net1492), .cc(net1457));
SW0 switch2815 (.gate(net266), .cc(net525));
SW0 switch2816 (.gate(net1357), .cc(net188));
SW switch2817 (.gate(cp1), .cc1(net246), .cc2(net123));
SW1 switch2818 (.gate(dor6), .cc(net7));
SW0 switch2819 (.gate(\0/ADL0 ), .cc(adl0));
SW0 switch2820 (.gate(net440), .cc(net813));
SW0 switch2821 (.gate(net335), .cc(net1280));
SW0 switch2822 (.gate(a1), .cc(net1549));
SW0 switch2823 (.gate(\PD-xxx010x1 ), .cc(\~TWOCYCLE ));
SW switch2824 (.gate(cp1), .cc1(net1650), .cc2(net94));
SW switch2825 (.gate(cclk), .cc1(net1602), .cc2(net506));
SW0 switch2826 (.gate(\notRdy0.delay ), .cc(net853));
SW0 switch2827 (.gate(net249), .cc(net163));
SW0 switch2828 (.gate(net249), .cc(dpc34_PCLC));
SW0 switch2829 (.gate(x2), .cc(notx2));
SW0 switch2830 (.gate(ir5), .cc(\op-sty/cpy-mem ));
SW0 switch2831 (.gate(ir5), .cc(\op-T0-iny/dey ));
SW0 switch2832 (.gate(ir5), .cc(\x-op-T0-tya ));
SW0 switch2833 (.gate(ir5), .cc(\op-T0-cpy/iny ));
SW0 switch2834 (.gate(ir5), .cc(\x-op-T0-txa ));
SW0 switch2835 (.gate(ir5), .cc(\op-T0-dex ));
SW0 switch2836 (.gate(ir5), .cc(\op-from-x ));
SW0 switch2837 (.gate(ir5), .cc(\op-T0-txs ));
SW0 switch2838 (.gate(ir5), .cc(\op-T+-dex ));
SW0 switch2839 (.gate(ir5), .cc(\op-T+-iny/dey ));
SW0 switch2840 (.gate(ir5), .cc(\op-T5-brk ));
SW0 switch2841 (.gate(ir5), .cc(\op-T0-php/pha ));
SW0 switch2842 (.gate(ir5), .cc(\op-T5-rti ));
SW0 switch2843 (.gate(ir5), .cc(\op-T0-eor ));
SW0 switch2844 (.gate(ir5), .cc(\op-T0-ora ));
SW0 switch2845 (.gate(ir5), .cc(\op-T4-rti ));
SW0 switch2846 (.gate(ir5), .cc(\op-T0-cmp ));
SW0 switch2847 (.gate(ir5), .cc(\op-T0-tya ));
SW0 switch2848 (.gate(ir5), .cc(\op-T0-txa ));
SW0 switch2849 (.gate(ir5), .cc(\op-T2-pha ));
SW0 switch2850 (.gate(ir5), .cc(\op-T2-brk ));
SW0 switch2851 (.gate(ir5), .cc(\op-sta/cmp ));
SW0 switch2852 (.gate(ir5), .cc(\op-T0-brk/rti ));
SW0 switch2853 (.gate(ir5), .cc(\op-brk/rti ));
SW0 switch2854 (.gate(ir5), .cc(\op-store ));
SW0 switch2855 (.gate(ir5), .cc(\op-T4-brk ));
SW0 switch2856 (.gate(ir5), .cc(\op-T2-php ));
SW0 switch2857 (.gate(ir5), .cc(\op-T2-php/pha ));
SW0 switch2858 (.gate(ir5), .cc(\op-T2-jmp-abs ));
SW0 switch2859 (.gate(ir5), .cc(\x-op-T4-rti ));
SW0 switch2860 (.gate(ir5), .cc(\op-T+-cmp ));
SW0 switch2861 (.gate(pipeUNK09), .cc(net941));
SW0 switch2862 (.gate(net256), .cc(net25));
SW switch2863 (.gate(cclk), .cc1(net633), .cc2(net1059));
SW switch2864 (.gate(cclk), .cc1(net1575), .cc2(pipeT2out));
SW0 switch2865 (.gate(net61), .cc(net1554));
SW0 switch2866 (.gate(net61), .cc(net479));
SW0 switch2867 (.gate(x4), .cc(notx4));
SW0 switch2868 (.gate(net479), .cc(dasb6));
SW0 switch2869 (.gate(notdor4), .cc(dor4));
SW0 switch2870 (.gate(\op-jsr ), .cc(net134));
SW0 switch2871 (.gate(notdor3), .cc(dor3));
SW0 switch2872 (.gate(\~op-branch-bit6 ), .cc(net1433));
SW1 switch2873 (.gate(net1315), .cc(net381));
SW switch2874 (.gate(net83), .cc1(net949), .cc2(net523));
SW0 switch2875 (.gate(net83), .cc(net1406));
SW0 switch2876 (.gate(AxB5), .cc(net570));
SW switch2877 (.gate(cclk), .cc1(net799), .cc2(\~NMIG ));
SW switch2878 (.gate(cclk), .cc1(net1693), .cc2(\~NMIG ));
SW0 switch2879 (.gate(net992), .cc(net46));
SW0 switch2880 (.gate(\op-T+-cmp ), .cc(\~op-set-C ));
SW0 switch2881 (.gate(net745), .cc(net241));
SW0 switch2882 (.gate(\branch-back.phi1 ), .cc(net1446));
SW switch2883 (.gate(\branch-back.phi1 ), .cc1(\short-circuit-branch-add ), .cc2(\~~alucout ));
SW switch2884 (.gate(net1184), .cc1(net474), .cc2(net766));
SW0 switch2885 (.gate(net1184), .cc(net410));
SW0 switch2886 (.gate(clearIR), .cc(\pd2.clearIR ));
SW0 switch2887 (.gate(clearIR), .cc(\pd6.clearIR ));
SW0 switch2888 (.gate(net838), .cc(net811));
SW0 switch2889 (.gate(ir4), .cc(notir4));
SW0 switch2890 (.gate(\~pchp1 ), .cc(pchp1));
SW switch2891 (.gate(cp1), .cc1(notRnWprepad), .cc2(net759));
SW0 switch2892 (.gate(idb0), .cc(net1687));
SW0 switch2893 (.gate(cclk), .cc(\~DBE ));
SW0 switch2894 (.gate(net541), .cc(ir7));
SW switch2895 (.gate(dpc20_ADDSB06), .cc1(alu1), .cc2(sb1));
SW0 switch2896 (.gate(pipeUNK12), .cc(net587));
SW switch2897 (.gate(dpc20_ADDSB06), .cc1(alu0), .cc2(dasb0));
SW0 switch2898 (.gate(net902), .cc(net1109));
SW0 switch2899 (.gate(net902), .cc(net1109));
SW0 switch2900 (.gate(net902), .cc(net1289));
SW0 switch2901 (.gate(net830), .cc(net1047));
SW1 switch2902 (.gate(net830), .cc(dpc23_SBAC));
SW0 switch2903 (.gate(net1643), .cc(net766));
SW0 switch2904 (.gate(net1643), .cc(dpc34_PCLC));
SW0 switch2905 (.gate(net1643), .cc(net410));
SW0 switch2906 (.gate(clearIR), .cc(\pd3.clearIR ));
SW0 switch2907 (.gate(clearIR), .cc(\pd4.clearIR ));
SW switch2908 (.gate(net1044), .cc1(net1408), .cc2(net1000));
SW switch2909 (.gate(cclk), .cc1(net1379), .cc2(pipeUNK10));
SW switch2910 (.gate(net986), .cc1(net1279), .cc2(net345));
SW switch2911 (.gate(dpc33_PCHDB), .cc1(pchp0), .cc2(idb0));
SW switch2912 (.gate(dpc33_PCHDB), .cc1(idb1), .cc2(pchp1));
SW switch2913 (.gate(dpc33_PCHDB), .cc1(idb2), .cc2(pchp2));
SW switch2914 (.gate(dpc33_PCHDB), .cc1(pchp3), .cc2(idb3));
SW switch2915 (.gate(dpc33_PCHDB), .cc1(pchp4), .cc2(idb4));
SW switch2916 (.gate(dpc33_PCHDB), .cc1(pchp5), .cc2(idb5));
SW switch2917 (.gate(dpc33_PCHDB), .cc1(idb6), .cc2(pchp6));
SW switch2918 (.gate(dpc33_PCHDB), .cc1(idb7), .cc2(pchp7));
SW switch2919 (.gate(cclk), .cc1(\~ABH5 ), .cc2(net869));
SW0 switch2920 (.gate(net1674), .cc(net772));
SW0 switch2921 (.gate(t5), .cc(\op-T5-rti/rts ));
SW0 switch2922 (.gate(t5), .cc(\xx-op-T5-jsr ));
SW0 switch2923 (.gate(t5), .cc(\op-T5-rts ));
SW0 switch2924 (.gate(t5), .cc(\op-T5-ind-x ));
SW0 switch2925 (.gate(t5), .cc(\op-T5-mem-ind-idx ));
SW0 switch2926 (.gate(t5), .cc(\op-T5-brk ));
SW0 switch2927 (.gate(t5), .cc(\op-T5-rti ));
SW0 switch2928 (.gate(t5), .cc(\op-T5-jsr ));
SW0 switch2929 (.gate(t5), .cc(\op-T5-ind-y ));
SW switch2930 (.gate(cclk), .cc1(net104), .cc2(net1221));
SW0 switch2931 (.gate(cclk), .cc(dpc3_SBX));
SW0 switch2932 (.gate(cclk), .cc(dpc2_XSB));
SW0 switch2933 (.gate(cclk), .cc(dpc1_SBY));
SW0 switch2934 (.gate(cclk), .cc(dpc0_YSB));
SW switch2935 (.gate(cp1), .cc1(net47), .cc2(net420));
SW0 switch2936 (.gate(net937), .cc(net1706));
SW0 switch2937 (.gate(net937), .cc(dpc34_PCLC));
SW0 switch2938 (.gate(net937), .cc(net1345));
SW0 switch2939 (.gate(net1132), .cc(net717));
SW switch2940 (.gate(cp1), .cc1(net666), .cc2(net1380));
SW0 switch2941 (.gate(\brk-done ), .cc(net334));
SW1 switch2942 (.gate(net617), .cc(net676));
SW switch2943 (.gate(cp1), .cc1(net1474), .cc2(notdor1));
SW0 switch2944 (.gate(net630), .cc(net1705));
SW0 switch2945 (.gate(net1518), .cc(dpc39_PCLPCL));
SW0 switch2946 (.gate(irline3), .cc(\op-T+-cpx/cpy-imm/zp ));
SW0 switch2947 (.gate(irline3), .cc(\op-sty/cpy-mem ));
SW0 switch2948 (.gate(irline3), .cc(\op-T0-iny/dey ));
SW0 switch2949 (.gate(irline3), .cc(\x-op-T0-tya ));
SW0 switch2950 (.gate(irline3), .cc(\op-T0-cpy/iny ));
SW0 switch2951 (.gate(irline3), .cc(\op-T0-cpx/inx ));
SW0 switch2952 (.gate(irline3), .cc(\op-T+-inx ));
SW0 switch2953 (.gate(irline3), .cc(\op-T+-iny/dey ));
SW0 switch2954 (.gate(irline3), .cc(\op-T0-ldy-mem ));
SW0 switch2955 (.gate(irline3), .cc(\op-T0-tay/ldy-not-idx ));
SW0 switch2956 (.gate(irline3), .cc(\op-T0-jsr ));
SW0 switch2957 (.gate(irline3), .cc(\op-T5-brk ));
SW0 switch2958 (.gate(irline3), .cc(\op-T0-php/pha ));
SW0 switch2959 (.gate(irline3), .cc(\op-T4-rts ));
SW0 switch2960 (.gate(irline3), .cc(\op-T3-plp/pla ));
SW0 switch2961 (.gate(irline3), .cc(\op-T5-rti ));
SW0 switch2962 (.gate(irline3), .cc(\op-jmp ));
SW0 switch2963 (.gate(irline3), .cc(\op-T2-stack ));
SW0 switch2964 (.gate(irline3), .cc(\op-T3-stack/bit/jmp ));
SW0 switch2965 (.gate(irline3), .cc(\op-T4-brk/jsr ));
SW0 switch2966 (.gate(irline3), .cc(\op-T4-rti ));
SW0 switch2967 (.gate(irline3), .cc(\op-plp/pla ));
SW0 switch2968 (.gate(irline3), .cc(\op-rti/rts ));
SW0 switch2969 (.gate(irline3), .cc(\op-T2-jsr ));
SW0 switch2970 (.gate(irline3), .cc(\op-T0-cpx/cpy/inx/iny ));
SW0 switch2971 (.gate(irline3), .cc(\op-T3-jmp ));
SW0 switch2972 (.gate(irline3), .cc(\op-T5-jsr ));
SW0 switch2973 (.gate(irline3), .cc(\op-T2-stack-access ));
SW0 switch2974 (.gate(irline3), .cc(\op-T0-tya ));
SW0 switch2975 (.gate(irline3), .cc(\op-T0-pla ));
SW0 switch2976 (.gate(irline3), .cc(\op-T0-tay ));
SW0 switch2977 (.gate(irline3), .cc(\op-T0-bit ));
SW0 switch2978 (.gate(irline3), .cc(\op-branch-done ));
SW0 switch2979 (.gate(irline3), .cc(\op-T2-pha ));
SW0 switch2980 (.gate(irline3), .cc(\op-T2-brk ));
SW0 switch2981 (.gate(irline3), .cc(\op-T3-jsr ));
SW0 switch2982 (.gate(irline3), .cc(\op-T2-branch ));
SW0 switch2983 (.gate(irline3), .cc(\op-T5-rts ));
SW0 switch2984 (.gate(irline3), .cc(\op-T0-brk/rti ));
SW0 switch2985 (.gate(irline3), .cc(\op-T0-jmp ));
SW0 switch2986 (.gate(irline3), .cc(\op-T3-branch ));
SW0 switch2987 (.gate(irline3), .cc(\op-brk/rti ));
SW0 switch2988 (.gate(irline3), .cc(\op-jsr ));
SW0 switch2989 (.gate(irline3), .cc(\x-op-jmp ));
SW0 switch2990 (.gate(irline3), .cc(\op-push/pull ));
SW0 switch2991 (.gate(irline3), .cc(\op-T4-brk ));
SW0 switch2992 (.gate(irline3), .cc(\op-T2-php ));
SW0 switch2993 (.gate(irline3), .cc(\op-T2-php/pha ));
SW0 switch2994 (.gate(irline3), .cc(\op-T4-jmp ));
SW0 switch2995 (.gate(irline3), .cc(\op-T5-rti/rts ));
SW0 switch2996 (.gate(irline3), .cc(\xx-op-T5-jsr ));
SW0 switch2997 (.gate(irline3), .cc(\op-T2-jmp-abs ));
SW0 switch2998 (.gate(irline3), .cc(\x-op-T3-plp/pla ));
SW0 switch2999 (.gate(irline3), .cc(\op-T0-cli/sei ));
SW0 switch3000 (.gate(irline3), .cc(\op-T+-bit ));
SW0 switch3001 (.gate(irline3), .cc(\op-T0-clc/sec ));
SW0 switch3002 (.gate(irline3), .cc(\x-op-T0-bit ));
SW0 switch3003 (.gate(irline3), .cc(\op-T0-plp ));
SW0 switch3004 (.gate(irline3), .cc(\x-op-T4-rti ));
SW0 switch3005 (.gate(irline3), .cc(\op-T+-cpx/cpy-abs ));
SW0 switch3006 (.gate(irline3), .cc(\x-op-push/pull ));
SW0 switch3007 (.gate(irline3), .cc(\op-T0-cld/sed ));
SW0 switch3008 (.gate(irline3), .cc(\op-clv ));
SW0 switch3009 (.gate(net312), .cc(net995));
SW switch3010 (.gate(net312), .cc1(net854), .cc2(net742));
SW0 switch3011 (.gate(net988), .cc(\~C34 ));
SW switch3012 (.gate(cp1), .cc1(net1291), .cc2(\brk-done ));
SW0 switch3013 (.gate(net717), .cc(RESG));
SW0 switch3014 (.gate(net717), .cc(net1087));
SW0 switch3015 (.gate(net1034), .cc(net1545));
SW1 switch3016 (.gate(net1034), .cc(net994));
SW0 switch3017 (.gate(pd7), .cc(\pd7.clearIR ));
SW0 switch3018 (.gate(idb3), .cc(DBZ));
SW0 switch3019 (.gate(pipeT2out), .cc(net1558));
SW0 switch3020 (.gate(pipeT2out), .cc(net12));
SW0 switch3021 (.gate(adl1), .cc(net1016));
SW0 switch3022 (.gate(net393), .cc(net551));
SW switch3023 (.gate(cclk), .cc1(pipeUNK23), .cc2(net1085));
SW switch3024 (.gate(cclk), .cc1(net1175), .cc2(pipeUNK28));
SW0 switch3025 (.gate(net1291), .cc(net1312));
SW switch3026 (.gate(\~C67 ), .cc1(net1013), .cc2(\~(AxBxC)7 ));
SW0 switch3027 (.gate(\~C67 ), .cc(\~(AxB7).C67 ));
SW0 switch3028 (.gate(\A+B1 ), .cc(net1510));
SW0 switch3029 (.gate(\pd1.clearIR ), .cc(\PD-0xx0xx0x ));
SW0 switch3030 (.gate(net90), .cc(Pout6));
SW0 switch3031 (.gate(net852), .cc(net1454));
SW0 switch3032 (.gate(net852), .cc(net260));
SW switch3033 (.gate(\op-inc/nop ), .cc1(net1107), .cc2(net1555));
SW0 switch3034 (.gate(net769), .cc(net1325));
SW1 switch3035 (.gate(net769), .cc(net1072));
SW0 switch3036 (.gate(pcl4), .cc(net1643));
SW switch3037 (.gate(net147), .cc1(db4), .cc2(db4));
SW0 switch3038 (.gate(net147), .cc(db4));
SW0 switch3039 (.gate(net147), .cc(db4));
SW0 switch3040 (.gate(net147), .cc(db4));
SW0 switch3041 (.gate(net147), .cc(db4));
SW0 switch3042 (.gate(net147), .cc(db4));
SW0 switch3043 (.gate(net147), .cc(db4));
SW0 switch3044 (.gate(net147), .cc(db4));
SW0 switch3045 (.gate(net147), .cc(db4));
SW0 switch3046 (.gate(idb2), .cc(net1376));
SW0 switch3047 (.gate(\PD-0xx0xx0x ), .cc(\PD-n-0xx0xx0x ));
SW0 switch3048 (.gate(\pipeT-SYNC ), .cc(net363));
SW0 switch3049 (.gate(net993), .cc(\~pclp6 ));
SW switch3050 (.gate(net753), .cc1(dasb5), .cc2(net1203));
SW0 switch3051 (.gate(net753), .cc(net1629));
SW0 switch3052 (.gate(RESG), .cc(D1x1));
SW switch3053 (.gate(cclk), .cc1(net632), .cc2(net339));
SW0 switch3054 (.gate(net1364), .cc(net108));
SW1 switch3055 (.gate(net1364), .cc(dpc16_EORS));
SW0 switch3056 (.gate(AxB1), .cc(\~(AxB)1 ));
SW0 switch3057 (.gate(net1467), .cc(cclk));
SW0 switch3058 (.gate(net1467), .cc(cclk));
SW0 switch3059 (.gate(net1467), .cc(cclk));
SW0 switch3060 (.gate(net1467), .cc(cclk));
SW0 switch3061 (.gate(pipeUNK34), .cc(net720));
SW0 switch3062 (.gate(net260), .cc(dasb7));
SW0 switch3063 (.gate(net735), .cc(dasb1));
SW0 switch3064 (.gate(adl2), .cc(net935));
SW0 switch3065 (.gate(net5), .cc(net146));
SW0 switch3066 (.gate(net1462), .cc(dpc38_PCLADL));
SW0 switch3067 (.gate(net1115), .cc(BRtaken));
SW0 switch3068 (.gate(notir5), .cc(\op-T0-cpx/inx ));
SW0 switch3069 (.gate(notir5), .cc(\op-T0-ldx/tax/tsx ));
SW0 switch3070 (.gate(notir5), .cc(\op-T+-inx ));
SW0 switch3071 (.gate(notir5), .cc(\op-T0-tsx ));
SW0 switch3072 (.gate(notir5), .cc(\op-T0-ldy-mem ));
SW0 switch3073 (.gate(notir5), .cc(\op-T0-tay/ldy-not-idx ));
SW0 switch3074 (.gate(notir5), .cc(\op-T0-jsr ));
SW0 switch3075 (.gate(notir5), .cc(\op-T4-rts ));
SW0 switch3076 (.gate(notir5), .cc(\op-T3-plp/pla ));
SW0 switch3077 (.gate(notir5), .cc(\op-ror ));
SW0 switch3078 (.gate(notir5), .cc(\op-plp/pla ));
SW0 switch3079 (.gate(notir5), .cc(\op-inc/nop ));
SW0 switch3080 (.gate(notir5), .cc(\op-T2-jsr ));
SW0 switch3081 (.gate(notir5), .cc(\op-T0-sbc ));
SW0 switch3082 (.gate(notir5), .cc(\op-T0-adc/sbc ));
SW0 switch3083 (.gate(notir5), .cc(\op-rol/ror ));
SW0 switch3084 (.gate(notir5), .cc(\op-T5-jsr ));
SW0 switch3085 (.gate(notir5), .cc(\op-T+-adc/sbc ));
SW0 switch3086 (.gate(notir5), .cc(\op-T0-pla ));
SW0 switch3087 (.gate(notir5), .cc(\op-T0-lda ));
SW0 switch3088 (.gate(notir5), .cc(\op-T0-tay ));
SW0 switch3089 (.gate(notir5), .cc(\op-T0-tax ));
SW0 switch3090 (.gate(notir5), .cc(\op-T0-bit ));
SW0 switch3091 (.gate(notir5), .cc(\op-T0-and ));
SW0 switch3092 (.gate(notir5), .cc(\op-T3-jsr ));
SW0 switch3093 (.gate(notir5), .cc(\op-T5-rts ));
SW0 switch3094 (.gate(notir5), .cc(\op-jsr ));
SW0 switch3095 (.gate(notir5), .cc(\xx-op-T5-jsr ));
SW0 switch3096 (.gate(notir5), .cc(\x-op-T3-plp/pla ));
SW0 switch3097 (.gate(notir5), .cc(\op-T+-bit ));
SW0 switch3098 (.gate(notir5), .cc(\x-op-T+-adc/sbc ));
SW0 switch3099 (.gate(notir5), .cc(\x-op-T0-bit ));
SW0 switch3100 (.gate(notir5), .cc(\op-T0-plp ));
SW0 switch3101 (.gate(notir5), .cc(\op-clv ));
SW0 switch3102 (.gate(pipeUNK41), .cc(net1497));
SW0 switch3103 (.gate(net1254), .cc(ab6));
SW0 switch3104 (.gate(net1254), .cc(ab6));
SW0 switch3105 (.gate(net1254), .cc(ab6));
SW0 switch3106 (.gate(net1254), .cc(ab6));
SW0 switch3107 (.gate(\pd4.clearIR ), .cc(\PD-xxx010x1 ));
SW0 switch3108 (.gate(\pd4.clearIR ), .cc(\PD-0xx0xx0x ));
SW0 switch3109 (.gate(\pd4.clearIR ), .cc(\PD-1xx000x0 ));
SW0 switch3110 (.gate(net236), .cc(net506));
SW0 switch3111 (.gate(net1580), .cc(net1656));
SW0 switch3112 (.gate(net1580), .cc(net1159));
SW switch3113 (.gate(net1573), .cc1(net845), .cc2(net1550));
SW0 switch3114 (.gate(\short-circuit-branch-add ), .cc(net959));
SW switch3115 (.gate(dpc2_XSB), .cc1(net578), .cc2(sb5));
SW switch3116 (.gate(dpc2_XSB), .cc1(net1724), .cc2(sb6));
SW0 switch3117 (.gate(net1256), .cc(dpc15_ANDS));
SW switch3118 (.gate(dpc2_XSB), .cc1(net1694), .cc2(sb2));
SW switch3119 (.gate(dpc2_XSB), .cc1(net242), .cc2(sb3));
SW switch3120 (.gate(dpc2_XSB), .cc1(net436), .cc2(dasb4));
SW0 switch3121 (.gate(net224), .cc(net520));
SW1 switch3122 (.gate(net224), .cc(net37));
SW0 switch3123 (.gate(net1719), .cc(net831));
SW0 switch3124 (.gate(\DA-C45 ), .cc(net570));
SW0 switch3125 (.gate(ir5), .cc(notir5));
SW0 switch3126 (.gate(notRdy0), .cc(fetch));
SW0 switch3127 (.gate(net1599), .cc(net538));
SW1 switch3128 (.gate(net1296), .cc(ab11));
SW0 switch3129 (.gate(irq), .cc(net1599));
SW switch3130 (.gate(cclk), .cc1(net1391), .cc2(pipeUNK15));
SW0 switch3131 (.gate(net531), .cc(net1255));
SW1 switch3132 (.gate(net531), .cc(dpc13_ORS));
SW1 switch3133 (.gate(dor7), .cc(net298));
SW switch3134 (.gate(cclk), .cc1(\~ABH4 ), .cc2(net999));
SW switch3135 (.gate(\ADH/ABH ), .cc1(net1298), .cc2(\~ABH1 ));
SW switch3136 (.gate(cclk), .cc1(net1106), .cc2(net1404));
SW0 switch3137 (.gate(notidl5), .cc(idl5));
SW0 switch3138 (.gate(notidl5), .cc(idl5));
SW0 switch3139 (.gate(notidl5), .cc(idl5));
SW0 switch3140 (.gate(\op-T4-rts ), .cc(net1464));
SW0 switch3141 (.gate(\op-T2-jsr ), .cc(net1649));
SW switch3142 (.gate(dpc0_YSB), .cc1(net767), .cc2(sb1));
SW switch3143 (.gate(alub1), .cc1(\~A.B1 ), .cc2(net189));
SW0 switch3144 (.gate(alub1), .cc(\~(A+B)1 ));
SW0 switch3145 (.gate(net662), .cc(dpc3_SBX));
SW0 switch3146 (.gate(net469), .cc(\~pchp5 ));
SW0 switch3147 (.gate(abl4), .cc(net86));
SW0 switch3148 (.gate(abl4), .cc(net1676));
SW1 switch3149 (.gate(abl4), .cc(net634));
SW0 switch3150 (.gate(notx1), .cc(net1709));
SW0 switch3151 (.gate(nots2), .cc(net1389));
SW0 switch3152 (.gate(\~A.B2 ), .cc(\DA-AB2 ));
SW0 switch3153 (.gate(net130), .cc(\ADL/ABL ));
SW0 switch3154 (.gate(net275), .cc(net104));
SW switch3155 (.gate(\PD-xxxx10x0 ), .cc1(net1515), .cc2(\~TWOCYCLE ));
SW0 switch3156 (.gate(\PD-xxxx10x0 ), .cc(net231));
SW0 switch3157 (.gate(\~pclp6 ), .cc(pclp6));
SW0 switch3158 (.gate(notRdy0), .cc(net1120));
SW switch3159 (.gate(notRdy0), .cc1(net1039), .cc2(net2));
SW0 switch3160 (.gate(\x-op-T3-ind-y ), .cc(net300));
SW0 switch3161 (.gate(\~(A+B)7 ), .cc(\A+B7 ));
SW0 switch3162 (.gate(\~(A+B)7 ), .cc(AxB7));
SW0 switch3163 (.gate(net617), .cc(net1140));
SW0 switch3164 (.gate(net1527), .cc(net1295));
SW0 switch3165 (.gate(\PD-n-0xx0xx0x ), .cc(net1515));
SW0 switch3166 (.gate(net1625), .cc(net90));
SW0 switch3167 (.gate(\x-op-T0-bit ), .cc(net1379));
SW0 switch3168 (.gate(net1697), .cc(net275));
SW0 switch3169 (.gate(\op-T5-ind-y ), .cc(net595));
SW0 switch3170 (.gate(\~(A+B)0 ), .cc(\DA-C01 ));
SW0 switch3171 (.gate(net782), .cc(net1347));
SW0 switch3172 (.gate(net366), .cc(\op-SRS ));
SW switch3173 (.gate(dpc39_PCLPCL), .cc1(pcl5), .cc2(pclp5));
SW switch3174 (.gate(dpc39_PCLPCL), .cc1(pcl4), .cc2(pclp4));
SW switch3175 (.gate(dpc39_PCLPCL), .cc1(pcl7), .cc2(pclp7));
SW switch3176 (.gate(dpc39_PCLPCL), .cc1(pcl6), .cc2(pclp6));
SW switch3177 (.gate(dpc39_PCLPCL), .cc1(pcl1), .cc2(pclp1));
SW switch3178 (.gate(dpc39_PCLPCL), .cc1(pcl0), .cc2(pclp0));
SW switch3179 (.gate(dpc39_PCLPCL), .cc1(pcl3), .cc2(pclp3));
SW switch3180 (.gate(dpc39_PCLPCL), .cc1(pcl2), .cc2(pclp2));
SW switch3181 (.gate(dpc27_SBADH), .cc1(adh5), .cc2(sb5));
SW switch3182 (.gate(dpc5_SADL), .cc1(net618), .cc2(adl6));
SW0 switch3183 (.gate(adh5), .cc(net254));
SW0 switch3184 (.gate(\~A.B6 ), .cc(net1038));
SW switch3185 (.gate(net1542), .cc1(net515), .cc2(net1158));
SW0 switch3186 (.gate(net1542), .cc(net1253));
SW0 switch3187 (.gate(net1247), .cc(dpc12_0ADD));
SW0 switch3188 (.gate(notidl1), .cc(idl1));
SW0 switch3189 (.gate(notidl1), .cc(idl1));
SW0 switch3190 (.gate(notidl1), .cc(idl1));
SW0 switch3191 (.gate(net1253), .cc(net515));
SW0 switch3192 (.gate(\op-SRS ), .cc(net160));
SW0 switch3193 (.gate(net837), .cc(\op-EORS ));
SW0 switch3194 (.gate(net590), .cc(alucin));
SW switch3195 (.gate(dpc4_SSB), .cc1(net332), .cc2(dasb0));
SW0 switch3196 (.gate(idb7), .cc(net423));
SW switch3197 (.gate(cclk), .cc1(pipeUNK02), .cc2(net774));
SW switch3198 (.gate(cclk), .cc1(\op-SRS ), .cc2(net968));
SW switch3199 (.gate(cclk), .cc1(\op-SUMS ), .cc2(net415));
SW switch3200 (.gate(cclk), .cc1(net680), .cc2(net1688));
SW0 switch3201 (.gate(net1528), .cc(net106));
SW0 switch3202 (.gate(\op-T0-bit ), .cc(net669));
SW switch3203 (.gate(dpc10_ADLADD), .cc1(adl6), .cc2(alub6));
SW switch3204 (.gate(dpc10_ADLADD), .cc1(adl7), .cc2(alub7));
SW1 switch3205 (.gate(net1608), .cc(ab13));
SW switch3206 (.gate(dpc10_ADLADD), .cc1(adl1), .cc2(alub1));
SW switch3207 (.gate(dpc10_ADLADD), .cc1(adl4), .cc2(alub4));
SW switch3208 (.gate(dpc10_ADLADD), .cc1(alub5), .cc2(adl5));
SW switch3209 (.gate(cclk), .cc1(net1126), .cc2(VEC0));
SW switch3210 (.gate(dpc10_ADLADD), .cc1(adl3), .cc2(alub3));
SW switch3211 (.gate(cclk), .cc1(net19), .cc2(pipeUNK18));
SW0 switch3212 (.gate(\dpc22_~DSA ), .cc(net1179));
SW0 switch3213 (.gate(net930), .cc(net1286));
SW0 switch3214 (.gate(db0), .cc(net718));
SW switch3216 (.gate(cclk), .cc1(net1618), .cc2(a2));
SW0 switch3217 (.gate(db2), .cc(net111));
SW switch3218 (.gate(cclk), .cc1(\~aluresult7 ), .cc2(notalu7));
SW0 switch3219 (.gate(db3), .cc(net896));
SW0 switch3220 (.gate(net1002), .cc(net1211));
SW switch3221 (.gate(net1416), .cc1(net1470), .cc2(net299));
SW0 switch3222 (.gate(net952), .cc(net152));
SW0 switch3223 (.gate(net862), .cc(net272));
SW switch3224 (.gate(\op-T2-idx-x-xy ), .cc1(net1717), .cc2(net1351));
SW switch3225 (.gate(dpc2_XSB), .cc1(net1709), .cc2(sb1));
SW0 switch3226 (.gate(net669), .cc(\op-ANDS ));
SW switch3228 (.gate(cclk), .cc1(NMIL), .cc2(net1252));
SW0 switch3229 (.gate(alua6), .cc(net1483));
SW0 switch3230 (.gate(alua6), .cc(\~(A+B)6 ));
SW0 switch3231 (.gate(net936), .cc(net1707));
SW0 switch3232 (.gate(net936), .cc(net388));
SW switch3233 (.gate(cclk), .cc1(a4), .cc2(net1344));
SW0 switch3234 (.gate(pch2), .cc(net1265));
SW0 switch3235 (.gate(noty7), .cc(net1251));
SW0 switch3236 (.gate(net865), .cc(net420));
SW0 switch3237 (.gate(NMIP), .cc(net645));
SW0 switch3238 (.gate(ir2), .cc(\op-T3-ind-y ));
SW0 switch3239 (.gate(ir2), .cc(\op-T2-abs-y ));
SW0 switch3240 (.gate(ir2), .cc(\op-T0-iny/dey ));
SW0 switch3241 (.gate(ir2), .cc(\x-op-T0-tya ));
SW0 switch3242 (.gate(ir2), .cc(\op-T2-ind-x ));
SW0 switch3243 (.gate(ir2), .cc(\x-op-T0-txa ));
SW0 switch3244 (.gate(ir2), .cc(\op-T0-dex ));
SW0 switch3245 (.gate(ir2), .cc(\op-T0-txs ));
SW0 switch3246 (.gate(ir2), .cc(\op-T+-dex ));
SW0 switch3247 (.gate(ir2), .cc(\op-T+-inx ));
SW0 switch3248 (.gate(ir2), .cc(\op-T0-tsx ));
SW0 switch3249 (.gate(ir2), .cc(\op-T+-iny/dey ));
SW0 switch3250 (.gate(ir2), .cc(\op-T0-jsr ));
SW0 switch3251 (.gate(ir2), .cc(\op-T5-brk ));
SW0 switch3252 (.gate(ir2), .cc(\op-T0-php/pha ));
SW0 switch3253 (.gate(ir2), .cc(\op-T4-rts ));
SW0 switch3254 (.gate(ir2), .cc(\op-T3-plp/pla ));
SW0 switch3255 (.gate(ir2), .cc(\op-T5-rti ));
SW0 switch3256 (.gate(ir2), .cc(\op-T2-stack ));
SW0 switch3257 (.gate(ir2), .cc(\op-T4-brk/jsr ));
SW0 switch3258 (.gate(ir2), .cc(\op-T4-rti ));
SW0 switch3259 (.gate(ir2), .cc(\op-T3-ind-x ));
SW0 switch3260 (.gate(ir2), .cc(\op-T4-ind-y ));
SW0 switch3261 (.gate(ir2), .cc(\op-T2-ind-y ));
SW0 switch3262 (.gate(ir2), .cc(\op-plp/pla ));
SW0 switch3263 (.gate(ir2), .cc(\op-T4-ind-x ));
SW0 switch3264 (.gate(ir2), .cc(\x-op-T3-ind-y ));
SW0 switch3265 (.gate(ir2), .cc(\op-rti/rts ));
SW0 switch3266 (.gate(ir2), .cc(\op-T2-jsr ));
SW0 switch3267 (.gate(ir2), .cc(\op-T5-jsr ));
SW0 switch3268 (.gate(ir2), .cc(\op-T2-stack-access ));
SW0 switch3269 (.gate(ir2), .cc(\op-T0-tya ));
SW0 switch3270 (.gate(ir2), .cc(\op-T+-shift-a ));
SW0 switch3271 (.gate(ir2), .cc(\op-T0-txa ));
SW0 switch3272 (.gate(ir2), .cc(\op-T0-pla ));
SW0 switch3273 (.gate(ir2), .cc(\op-T0-tay ));
SW0 switch3274 (.gate(ir2), .cc(\op-T0-shift-a ));
SW0 switch3275 (.gate(ir2), .cc(\op-T0-tax ));
SW0 switch3276 (.gate(ir2), .cc(\op-T5-ind-y ));
SW0 switch3277 (.gate(ir2), .cc(\op-branch-done ));
SW0 switch3278 (.gate(ir2), .cc(\op-T2-pha ));
SW0 switch3279 (.gate(ir2), .cc(\op-T0-shift-right-a ));
SW0 switch3280 (.gate(ir2), .cc(\op-T2-brk ));
SW0 switch3281 (.gate(ir2), .cc(\op-T3-jsr ));
SW0 switch3282 (.gate(ir2), .cc(\op-T2-branch ));
SW0 switch3283 (.gate(ir2), .cc(\op-T2-ind ));
SW0 switch3284 (.gate(ir2), .cc(\op-T5-rts ));
SW0 switch3285 (.gate(ir2), .cc(\op-T0-brk/rti ));
SW0 switch3286 (.gate(ir2), .cc(\op-T5-ind-x ));
SW0 switch3287 (.gate(ir2), .cc(\x-op-T4-ind-y ));
SW0 switch3288 (.gate(ir2), .cc(\op-T3-branch ));
SW0 switch3289 (.gate(ir2), .cc(\op-brk/rti ));
SW0 switch3290 (.gate(ir2), .cc(\op-jsr ));
SW0 switch3291 (.gate(ir2), .cc(\op-push/pull ));
SW0 switch3292 (.gate(ir2), .cc(\op-T4-brk ));
SW0 switch3293 (.gate(ir2), .cc(\op-T2-php ));
SW0 switch3294 (.gate(ir2), .cc(\op-T2-php/pha ));
SW0 switch3295 (.gate(ir2), .cc(\op-T5-rti/rts ));
SW0 switch3296 (.gate(ir2), .cc(\xx-op-T5-jsr ));
SW0 switch3297 (.gate(ir2), .cc(\x-op-T3-plp/pla ));
SW0 switch3298 (.gate(ir2), .cc(\op-T0-cli/sei ));
SW0 switch3299 (.gate(ir2), .cc(\op-T0-clc/sec ));
SW0 switch3300 (.gate(ir2), .cc(\op-T0-plp ));
SW0 switch3301 (.gate(ir2), .cc(\x-op-T4-rti ));
SW0 switch3302 (.gate(ir2), .cc(\op-T+-asl/rol-a ));
SW0 switch3303 (.gate(ir2), .cc(\x-op-push/pull ));
SW0 switch3304 (.gate(ir2), .cc(\op-T0-cld/sed ));
SW0 switch3305 (.gate(ir2), .cc(\op-T5-mem-ind-idx ));
SW0 switch3306 (.gate(ir2), .cc(\op-clv ));
SW0 switch3307 (.gate(ir2), .cc(\op-implied ));
SW switch3308 (.gate(cclk), .cc1(net1712), .cc2(pipeVectorA2));
SW0 switch3309 (.gate(notx7), .cc(net871));
SW0 switch3310 (.gate(\op-T5-ind-x ), .cc(net726));
SW0 switch3311 (.gate(\op-T5-ind-x ), .cc(net256));
SW0 switch3312 (.gate(net1463), .cc(net1076));
SW1 switch3313 (.gate(net1463), .cc(net147));
SW0 switch3314 (.gate(s1), .cc(net1711));
SW0 switch3315 (.gate(\op-T0-tya ), .cc(net1455));
SW switch3316 (.gate(cclk), .cc1(y0), .cc2(net564));
SW switch3317 (.gate(cclk), .cc1(net659), .cc2(\~ABH7 ));
SW0 switch3318 (.gate(net1213), .cc(net1209));
SW0 switch3319 (.gate(net228), .cc(dpc30_ADHPCH));
SW0 switch3320 (.gate(net1224), .cc(net186));
SW0 switch3321 (.gate(notalu3), .cc(alu3));
SW0 switch3322 (.gate(net1277), .cc(net1441));
SW1 switch3323 (.gate(net1277), .cc(\dpc42_DL/ADH ));
SW0 switch3324 (.gate(notRdy0), .cc(net781));
SW0 switch3325 (.gate(notRdy0), .cc(net781));
SW0 switch3326 (.gate(net134), .cc(net930));
SW0 switch3327 (.gate(net134), .cc(net467));
SW switch3328 (.gate(cclk), .cc1(pipephi2Reset0), .cc2(RESP));
SW0 switch3329 (.gate(net811), .cc(net1080));
SW switch3330 (.gate(net811), .cc1(net1205), .cc2(net100));
SW1 switch3331 (.gate(cclk), .cc(idb1));
SW0 switch3332 (.gate(\pd1.clearIR ), .cc(net1641));
SW switch3333 (.gate(net609), .cc1(net1192), .cc2(net1547));
SW switch3334 (.gate(net609), .cc1(net1209), .cc2(net1264));
SW0 switch3335 (.gate(net1412), .cc(net384));
SW0 switch3336 (.gate(db7), .cc(net62));
SW switch3337 (.gate(cp1), .cc1(net1338), .cc2(net720));
SW0 switch3338 (.gate(net1464), .cc(net1109));
SW switch3339 (.gate(cp1), .cc1(net227), .cc2(net703));
SW1 switch3340 (.gate(cclk), .cc(sb5));
SW switch3341 (.gate(cclk), .cc1(net548), .cc2(nots7));
SW switch3342 (.gate(cp1), .cc1(net1095), .cc2(idl4));
SW0 switch3343 (.gate(cp1), .cc(net43));
SW0 switch3344 (.gate(cp1), .cc(net839));
SW0 switch3345 (.gate(net1049), .cc(net507));
SW0 switch3346 (.gate(pipeUNK08), .cc(net954));
SW switch3347 (.gate(dpc11_SBADD), .cc1(sb7), .cc2(alua7));
SW0 switch3348 (.gate(y5), .cc(noty5));
SW0 switch3349 (.gate(net598), .cc(net1260));
SW0 switch3350 (.gate(net310), .cc(ir0));
SW0 switch3351 (.gate(adh7), .cc(net494));
SW1 switch3352 (.gate(cclk), .cc(adh6));
SW1 switch3353 (.gate(cclk), .cc(adl7));
SW0 switch3354 (.gate(net180), .cc(net501));
SW0 switch3355 (.gate(\~pclp1 ), .cc(pclp1));
SW switch3356 (.gate(\~op-branch-done ), .cc1(net239), .cc2(net192));
SW0 switch3357 (.gate(noty3), .cc(net1531));
SW switch3358 (.gate(cclk), .cc1(net1199), .cc2(notidl2));
SW switch3359 (.gate(cclk), .cc1(net824), .cc2(pipeUNK34));
SW0 switch3360 (.gate(cclk), .cc(net886));
SW switch3361 (.gate(\ADL/ABL ), .cc1(net524), .cc2(\~ABL6 ));
SW switch3362 (.gate(\ADL/ABL ), .cc1(net577), .cc2(\~ABL7 ));
SW switch3363 (.gate(\ADL/ABL ), .cc1(net738), .cc2(\~ABL4 ));
SW switch3364 (.gate(\ADL/ABL ), .cc1(net463), .cc2(\~ABL5 ));
SW0 switch3365 (.gate(adl5), .cc(net1094));
SW0 switch3366 (.gate(\~NMIG ), .cc(net1712));
SW0 switch3367 (.gate(\x-op-T4-ind-y ), .cc(net261));
SW0 switch3368 (.gate(\x-op-T4-ind-y ), .cc(net726));
SW switch3369 (.gate(fetch), .cc1(net380), .cc2(clearIR));
SW0 switch3370 (.gate(pipeUNK35), .cc(net238));
SW switch3371 (.gate(\~A.B0 ), .cc1(\DA-C01 ), .cc2(net1354));
SW0 switch3372 (.gate(\~ABH1 ), .cc(abh1));
SW switch3373 (.gate(dpc40_ADLPCL), .cc1(pcl1), .cc2(adl1));
SW switch3374 (.gate(dpc40_ADLPCL), .cc1(adl0), .cc2(pcl0));
SW switch3375 (.gate(dpc40_ADLPCL), .cc1(pcl3), .cc2(adl3));
SW switch3376 (.gate(dpc40_ADLPCL), .cc1(adl2), .cc2(pcl2));
SW switch3377 (.gate(dpc40_ADLPCL), .cc1(pcl5), .cc2(adl5));
SW switch3378 (.gate(dpc40_ADLPCL), .cc1(adl4), .cc2(pcl4));
SW switch3379 (.gate(dpc40_ADLPCL), .cc1(adl6), .cc2(pcl6));
SW0 switch3380 (.gate(notRdy0), .cc(\short-circuit-idx-add ));
SW0 switch3381 (.gate(idb0), .cc(DBZ));
SW0 switch3382 (.gate(net1271), .cc(dpc27_SBADH));
SW0 switch3383 (.gate(res), .cc(net312));
SW switch3384 (.gate(dpc20_ADDSB06), .cc1(alu2), .cc2(sb2));
SW0 switch3385 (.gate(net499), .cc(net1659));
SW0 switch3386 (.gate(net499), .cc(net743));
SW0 switch3387 (.gate(\op-T+-cpx/cpy-abs ), .cc(\~op-set-C ));
SW0 switch3388 (.gate(nots6), .cc(net618));
SW switch3389 (.gate(cclk), .cc1(net1341), .cc2(net695));
SW1 switch3390 (.gate(net475), .cc(ab12));
SW switch3391 (.gate(dpc6_SBS), .cc1(s7), .cc2(sb7));
SW0 switch3392 (.gate(net642), .cc(ab2));
SW0 switch3393 (.gate(net642), .cc(ab2));
SW0 switch3394 (.gate(net642), .cc(ab2));
SW0 switch3395 (.gate(net642), .cc(ab2));
SW0 switch3396 (.gate(net1002), .cc(net152));
SW0 switch3397 (.gate(net572), .cc(net1407));
SW switch3398 (.gate(cclk), .cc1(pipeUNK17), .cc2(net334));
SW1 switch3399 (.gate(net1479), .cc(ab1));
SW1 switch3400 (.gate(net1479), .cc(ab1));
SW1 switch3401 (.gate(net1479), .cc(ab1));
SW1 switch3402 (.gate(net1479), .cc(ab1));
SW1 switch3403 (.gate(net1479), .cc(ab1));
SW0 switch3404 (.gate(x3), .cc(notx3));
SW0 switch3405 (.gate(net323), .cc(net14));
SW0 switch3406 (.gate(net355), .cc(net593));
SW1 switch3407 (.gate(net355), .cc(dpc4_SSB));
SW0 switch3408 (.gate(net392), .cc(net814));
SW0 switch3409 (.gate(net392), .cc(net557));
SW0 switch3410 (.gate(net794), .cc(db1));
SW0 switch3411 (.gate(net794), .cc(db1));
SW0 switch3412 (.gate(net794), .cc(db1));
SW0 switch3413 (.gate(net794), .cc(db1));
SW0 switch3414 (.gate(net794), .cc(db1));
SW0 switch3415 (.gate(net794), .cc(db1));
SW0 switch3416 (.gate(net794), .cc(db1));
SW switch3417 (.gate(cclk), .cc1(\x-op-T+-adc/sbc ), .cc2(pipeUNK03));
SW switch3418 (.gate(cclk), .cc1(net696), .cc2(net610));
SW0 switch3419 (.gate(alucout), .cc(net811));
SW0 switch3420 (.gate(notRdy0), .cc(net1440));
SW0 switch3421 (.gate(\~A.B1 ), .cc(net936));
SW0 switch3422 (.gate(dor7), .cc(net1501));
SW0 switch3423 (.gate(dor7), .cc(net23));
SW0 switch3424 (.gate(net1247), .cc(dpc0_YSB));
SW0 switch3425 (.gate(net43), .cc(net1230));
SW0 switch3426 (.gate(net122), .cc(net570));
SW0 switch3427 (.gate(\~(A+B)3 ), .cc(\A+B3 ));
SW0 switch3428 (.gate(\~(A+B)3 ), .cc(AxB3));
SW0 switch3429 (.gate(alua2), .cc(net452));
SW0 switch3430 (.gate(alua2), .cc(\~(A+B)2 ));
SW0 switch3431 (.gate(\op-SRS ), .cc(\op-SUMS ));
SW0 switch3432 (.gate(cclk), .cc(net1585));
SW0 switch3433 (.gate(net1270), .cc(net1518));
SW1 switch3434 (.gate(net1270), .cc(dpc39_PCLPCL));
SW0 switch3435 (.gate(sb3), .cc(net432));
SW0 switch3436 (.gate(sb3), .cc(net432));
SW0 switch3437 (.gate(net906), .cc(net714));
SW0 switch3438 (.gate(net906), .cc(dpc19_ADDSB7));
SW0 switch3439 (.gate(notx5), .cc(net578));
SW0 switch3440 (.gate(net1338), .cc(net462));
SW0 switch3441 (.gate(\brk-done ), .cc(INTG));
SW1 switch3442 (.gate(net7), .cc(db6));
SW1 switch3443 (.gate(net7), .cc(db6));
SW1 switch3444 (.gate(net7), .cc(db6));
SW0 switch3445 (.gate(net680), .cc(net1526));
SW switch3446 (.gate(cclk), .cc1(net629), .cc2(net760));
SW0 switch3447 (.gate(nnT2BR), .cc(net1427));
SW0 switch3448 (.gate(sb7), .cc(net852));
SW0 switch3449 (.gate(sb7), .cc(net852));
SW0 switch3450 (.gate(net138), .cc(ab3));
SW0 switch3451 (.gate(net138), .cc(ab3));
SW0 switch3452 (.gate(net138), .cc(ab3));
SW0 switch3453 (.gate(net138), .cc(ab3));
SW switch3454 (.gate(cclk), .cc1(net1649), .cc2(net1027));
SW0 switch3455 (.gate(RESG), .cc(notRnWprepad));
SW switch3456 (.gate(net638), .cc1(net1118), .cc2(net604));
SW0 switch3457 (.gate(net1358), .cc(net396));
SW1 switch3458 (.gate(net634), .cc(ab4));
SW1 switch3459 (.gate(net634), .cc(ab4));
SW1 switch3460 (.gate(net634), .cc(ab4));
SW1 switch3461 (.gate(net634), .cc(ab4));
SW1 switch3462 (.gate(net634), .cc(ab4));
SW switch3463 (.gate(net1542), .cc1(net1099), .cc2(net1568));
SW switch3464 (.gate(net1253), .cc1(net1184), .cc2(net1498));
SW0 switch3465 (.gate(net1253), .cc(net903));
SW0 switch3466 (.gate(D1x1), .cc(net1471));
SW0 switch3467 (.gate(net386), .cc(net392));
SW0 switch3468 (.gate(net386), .cc(dpc34_PCLC));
SW switch3469 (.gate(cclk), .cc1(net700), .cc2(net1565));
SW0 switch3470 (.gate(net329), .cc(net1166));
SW0 switch3471 (.gate(net329), .cc(dpc34_PCLC));
SW0 switch3472 (.gate(\op-T4-ind-y ), .cc(net1107));
SW0 switch3473 (.gate(net1072), .cc(db0));
SW0 switch3474 (.gate(net1072), .cc(db0));
SW0 switch3475 (.gate(net1072), .cc(db0));
SW0 switch3476 (.gate(net1072), .cc(db0));
SW0 switch3477 (.gate(net1072), .cc(db0));
SW0 switch3478 (.gate(net1072), .cc(db0));
SW0 switch3479 (.gate(net1072), .cc(db0));
SW0 switch3480 (.gate(net1072), .cc(db0));
SW switch3481 (.gate(\~C45 ), .cc1(\~(AxBxC)5 ), .cc2(net547));
SW0 switch3482 (.gate(\~C45 ), .cc(\~(AxB5).C45 ));
SW1 switch3483 (.gate(net826), .cc(ab8));
SW0 switch3484 (.gate(net218), .cc(net1716));
SW switch3485 (.gate(cclk), .cc1(net1594), .cc2(net688));
SW0 switch3486 (.gate(net1395), .cc(RESP));
SW0 switch3487 (.gate(net1395), .cc(RESP));
SW switch3488 (.gate(pipeUNK10), .cc1(net941), .cc2(net1111));
SW switch3489 (.gate(dpc13_ORS), .cc1(\~(A+B)1 ), .cc2(\~aluresult1 ));
SW0 switch3490 (.gate(\op-T0-and ), .cc(net669));
SW0 switch3491 (.gate(net6), .cc(net282));
SW1 switch3492 (.gate(net6), .cc(dpc6_SBS));
SW switch3493 (.gate(\op-sta/cmp ), .cc1(net1280), .cc2(net1037));
SW0 switch3494 (.gate(net43), .cc(net35));
SW0 switch3495 (.gate(idb1), .cc(net583));
SW0 switch3496 (.gate(x6), .cc(notx6));
SW0 switch3497 (.gate(net678), .cc(t3));
SW switch3498 (.gate(cclk), .cc1(pd1), .cc2(net1319));
SW switch3499 (.gate(cclk), .cc1(pd0), .cc2(net93));
SW0 switch3500 (.gate(net951), .cc(net1152));
SW1 switch3501 (.gate(net951), .cc(net642));
SW1 switch3502 (.gate(cclk), .cc(sb2));
SW switch3503 (.gate(cclk), .cc1(net1190), .cc2(nots2));
SW1 switch3504 (.gate(cclk), .cc(idb4));
SW0 switch3505 (.gate(net1258), .cc(net1130));
SW0 switch3506 (.gate(net1619), .cc(net586));
SW0 switch3507 (.gate(net923), .cc(net356));
SW0 switch3508 (.gate(net923), .cc(dpc35_PCHC));
SW0 switch3509 (.gate(net923), .cc(net810));

endmodule
