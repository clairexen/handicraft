module testbox_1(input A, B, output Y);
assign Y = 1;
endmodule
