module test011(a0, a1, a2, a3, y);
  wire [1:0] _00_;
  wire _01_;
  wire _02_;
  wire _03_;
  wire _04_;
  wire _05_;
  wire _06_;
  wire _07_;
  wire _08_;
  wire _09_;
  wire _10_;
  wire _11_;
  wire [4:0] _12_;
  wire [3:0] _13_;
  wire [3:0] _14_;
  input [3:0] a0;
  input [3:0] a1;
  input [3:0] a2;
  input [3:0] a3;
  output [44:0] y;
  wire [4:0] y1;
  wire [5:0] y2;
  wire [3:0] y3;
  wire [4:0] y4;
  wire [3:0] y5;
  assign _14_[0] = a0[0] ^ a1[0];
  assign _14_[1] = a0[1] ^ a1[1];
  assign _14_[2] = a0[2] ^ a1[2];
  assign _14_[3] = a0[3] ^ a1[3];
  assign _00_[0] = _14_[0] | _14_[1];
  assign _00_[1] = _14_[2] | _14_[3];
  assign y[40] = _00_[0] | _00_[1];
  assign y[30] = ~_12_[4];
  assign _13_[1] = ~a2[1];
  assign _13_[2] = ~a2[2];
  assign _13_[3] = ~a2[3];
  assign _13_[0] = ~a2[0];
  assign _01_ = a3[0] & _13_[0];
  assign _02_ = a3[0] ^ _13_[0];
  assign _12_[1] = _01_ | _02_;
  assign _03_ = a3[1] & _13_[1];
  assign _04_ = a3[1] ^ _13_[1];
  assign _05_ = _04_ & _12_[1];
  assign _12_[2] = _03_ | _05_;
  assign _06_ = a3[2] & _13_[2];
  assign _07_ = a3[2] ^ _13_[2];
  assign _08_ = _07_ & _12_[2];
  assign _12_[3] = _06_ | _08_;
  assign _09_ = a3[3] & _13_[3];
  assign _10_ = a3[3] ^ _13_[3];
  assign _11_ = _10_ & _12_[3];
  assign _12_[4] = _09_ | _11_;
  assign { y[44:41], y[39:31], y[29:0] } = { 6'b000000, a0, 7'b0000000, y[40], y[30], y[30], y[30], y[30], 21'b000000000000000000000 };
  assign y1 = { 4'b0000, y[40] };
  assign y2 = { 2'b00, a0 };
  assign y3 = { 3'b000, y[30] };
  assign y4 = { 4'b0000, y[40] };
  assign y5 = { y[30], y[30], y[30], y[30] };
endmodule
