module testbench;
	reg clk;
	always #5 clk = (clk === 1'b0);

	integer cycles = 0;

	always @(posedge clk)
		cycles <= cycles + 1;

	reg         pdep;
	reg         pext;
	reg  [63:0] din;
	reg  [63:0] mask;
	wire [63:0] dout;

`ifdef PDEP_PEXT_MC
	reg load;
	wire ready;

	pdep_pext_mc3 uut (
		.clk   (clk  ),
		.load  (load ),
		.pext  (pext ),
		.ready (ready),
		.din   (din  ),
		.mask  (mask ),
		.dout  (dout )
	);
`else
	pdep_pext uut (
		.pdep (pdep),
		.pext (pext),
		.din  (din ),
		.mask (mask),
		.dout (dout)
	);
`endif

	integer test_count = 0;

	task test (
		input [63:0] i_value,
		input [63:0] i_mask,
		input [63:0] o_pext,
		input [63:0] o_pdep,
		input [63:0] o_grev
	);
		begin
`ifdef PDEP_PEXT_MC
			din <= i_value;
			mask <= i_mask;
			pext <= 0;
			load <= 1;
			@(posedge clk);

			load <= 0;
			while (!ready) @(posedge clk);

			if (dout != o_pdep) begin
				$display("Error in PDEP!");
				$display("  value  = %x", din);
				$display("  mask   = %x", mask);
				$display("  result = %x", dout);
				$display("  expect = %x", o_pdep);
				@(posedge clk);
				@(posedge clk);
				$stop;
			end

			pext <= 1;
			load <= 1;
			@(posedge clk);

			load <= 0;
			while (!ready) @(posedge clk);

			if (dout != o_pext) begin
				$display("Error in PEXT!");
				$display("  value  = %x", din);
				$display("  mask   = %x", mask);
				$display("  result = %x", dout);
				$display("  expect = %x", o_pext);
				@(posedge clk);
				@(posedge clk);
				$stop;
			end
`else
			din <= i_value;
			mask <= i_mask;

			pdep <= 1;
			pext <= 0;
			@(posedge clk);

			if (dout != o_pdep) begin
				$display("Error in PDEP!");
				$display("  value  = %x", din);
				$display("  mask   = %x", mask);
				$display("  result = %x", dout);
				$display("  expect = %x", o_pdep);
				@(posedge clk);
				@(posedge clk);
				$stop;
			end

			pdep <= 0;
			pext <= 1;
			@(posedge clk);

			if (dout != o_pext) begin
				$display("Error in PEXT!");
				$display("  value  = %x", din);
				$display("  mask   = %x", mask);
				$display("  result = %x", dout);
				$display("  expect = %x", o_pext);
				@(posedge clk);
				@(posedge clk);
				$stop;
			end

			pdep <= 0;
			pext <= 0;
			@(posedge clk);

			if (dout != o_grev) begin
				$display("Error in GREV!");
				$display("  value  = %x", din);
				$display("  mask   = %x", mask);
				$display("  result = %x", dout);
				$display("  expect = %x", o_grev);
				@(posedge clk);
				@(posedge clk);
				$stop;
			end
`endif
			test_count = test_count + 1;
			if (test_count % 100 == 0) begin
				$display("Completed %1d tests.", test_count);
			end
		end
	endtask

	initial begin
		$dumpfile("testbench.vcd");
		$dumpvars(0, testbench);

		// generated by model.cc
		test(64'h79690975fbde15b0, 64'h2a337357ae2cc59b, 64'h00000003487bd678, 64'h0a3333170208c180, 64'hea0969e9d08ab7fd);
		test(64'h2fef107a27529ad0, 64'he4093df8432a8be5, 64'h000000001e87b3d8, 64'h4009292801220a80, 64'hb11a560ef1fd025b);
		test(64'h71dd0913271687b2, 64'hf70abb341875063d, 64'h00000000730a8378, 64'h2308131000350224, 64'h17b492b13260ee2b);
		test(64'h61b97bcd4b21c371, 64'he845105ed8c77cb7, 64'h00000000c7650c19, 64'ha004104408c034a1, 64'hc38ed284deb3869d);
		test(64'he77b20aec4233f8e, 64'hc9ddc8f042775a71, 64'h00000001ae8a9370, 64'h4810403000774070, 64'h3f4dc813105ddbb7);
		test(64'hfe5defe9c5610885, 64'h6ef14999f8114bd4, 64'h00000000fafde149, 64'h60a1400810004044, 64'hfe9eefd580585c16);
		test(64'ha3a03fe4de4f1c43, 64'h9fded21c82caf2bb, 64'h00000008e033b883, 64'h135c401c800a8203, 64'h2c832fb772cf505c);
		test(64'hb494d6880418a99e, 64'h955753b579933f4d, 64'h0000001cce801296, 64'h100010050882194c, 64'h8687449e4280d665);
		test(64'h01239ff2c4a06a73, 64'h8be87413a8b3d667, 64'h00000000247a613b, 64'h0a20240000a28643, 64'h230556ce80c4f94f);
		test(64'h2e6f66b049cdc80b, 64'hf991db0c819b315b, 64'h0000000028a43507, 64'h48118a0c80100013, 64'hd0666f470d313b29);
		test(64'h94269b57fb8d31f9, 64'hbe1edefcfabd75da, 64'h00000a8ed57f9dbe, 64'h9a0adeb8321835c2, 64'h5d6e8961f6c427fe);
		test(64'he35ac67471cc39b1, 64'h7b59baf2b613ed82, 64'h0000000cfa2e6036, 64'h215038601601a802, 64'hbc5a39d1d433c6e4);
		test(64'h8b4eb7817f86ead9, 64'h97876671a300714c, 64'h0000000009b38be6, 64'h9700626121005104, 64'he4b8187b68f79dae);
		test(64'hfad4dc52cb2fa2ae, 64'h11e69a347dd2966b, 64'h000000016b94a32e, 64'h018490247902122a, 64'h4f3d5754b2f5a4b3);
		test(64'h686f3326a04fc987, 64'h6ed5ff7aa865d7d4, 64'h000000e2ccd3af19, 64'h08c4811aa8045054, 64'h336286f69c780af4);
		test(64'h6edd22562c4c697b, 64'h5b22f45380f3cf69, 64'h00000001609c419f, 64'h0222101200624749, 64'h8c1cb796ee9da911);
		test(64'haf29109cc782d2b7, 64'h76d874a3714b9ad2, 64'h00000000b12892db, 64'h3058400261028a52, 64'h4063af8678ed3d28);
		test(64'h7dc2ae94e4dbf967, 64'h0c971bea6a6af755, 64'h0000000726865f9b, 64'h081608ca2a6a2615, 64'hd586eb1c6fb98d7e);
		test(64'hea2177d8d51f57fb, 64'h76104a9e26b7f794, 64'h0000000195e23d7e, 64'h320042062625f714, 64'h778dae1275bf5df1);
		test(64'h6d159abfb303fd7b, 64'h0ff20e6dfbb7c441, 64'h000000068abed87f, 64'h0f600c00fb93c041, 64'h9e2a657f7303feb7);
		test(64'hd251a40a022b9b89, 64'h6c129af7f2440efe, 64'h00000002280412c4, 64'h40000825c2400e12, 64'h62e6e880a01a4587);
		test(64'hc7dee68fffbaf963, 64'h15ada4e53975b451, 64'h0000000076f3f675, 64'h15ad84c43944a011, 64'hd94fcbedf693ff75);
		test(64'h63eb500cce126b79, 64'h314320aa7da5b1ef, 64'h00000000bc5302b9, 64'h3003200048a130e9, 64'h48739ed6d7c6300a);
		test(64'hd27d2fde3497614c, 64'hbe55668178139c8e, 64'h0000000053ef3706, 64'h3410468060011088, 64'h7d87b7f8d61c3149);
		test(64'h9480583abdfb5837, 64'h9d8dbb3a5bde4347, 64'h0000001a833dbec7, 64'h9485ab3852c00307, 64'h29011a5cbddf1aec);
		test(64'h61fd04828c93ce01, 64'hdf9a26c8470349dd, 64'h0000000043ca2781, 64'h861020c841030001, 64'h1480ef2920dc36c4);
		test(64'hca9d54bd4e78980e, 64'hb1db9b0fecbfaabe, 64'h00000116a356e287, 64'h21d28309e026001c, 64'hb0262db17e1576a3);
		test(64'he79541e25d0dba6b, 64'hff98837fda2a5bdf, 64'h000001cf8e27272b, 64'hf1080350ca0a48cb, 64'h4782a9e7d65db0ba);
		test(64'hc3bd5e2cd52318a8, 64'h02ab7bb54e687499, 64'h00000000f6e5522a, 64'h0289221406005080, 64'h1cad7ec3542413ea);
		test(64'hbebf0929f41aa230, 64'h58aee9fdc3f41b74, 64'h0000000fe32b8226, 64'h102ea01941100300, 64'h2a034fa19092ebfb);
		test(64'h62daff171a9fae42, 64'he5baa16ee5b5419e, 64'h000000032fc60b81, 64'he032202ec4b04004, 64'hd4ffa78981baf6a4);
		test(64'h16b3a918e4278c9d, 64'h4ab9cfc9a41744c4, 64'h000000000f692eed, 64'h40808780a0044484, 64'h613b9a814e72c8d9);
		test(64'h86ddce906c8cdb4d, 64'h867e3492977cb1bb, 64'h00000007b8e20ec5, 64'h003604009158a119, 64'h2bbd13639037bb16);
		test(64'h3d0e482377794618, 64'h90e1bc8ba22d3294, 64'h0000000004046f4a, 64'h10c1b08202201200, 64'h8432d3e064817797);
		test(64'hf48119b103954df1, 64'h79780d4e5b2b3b2a, 64'h00000001c0a0312c, 64'h4018084448293a02, 64'h650cf41724f1e446);
		test(64'hb36eb1caa58ee7dc, 64'hf0fe55be95a18d13, 64'h00000005b7596e5c, 64'h504a40b681a18510, 64'hd835dc677eb35a17);
		test(64'h1234769364d9eac9, 64'h31a7445bdf8bcb5c, 64'h0000000266b49bea, 64'h112440198f094844, 64'h396743219cae9d46);
		test(64'h1735808ee4398bca, 64'h8f09996552504a5d, 64'h0000000003b05174, 64'h0801906010504814, 64'hd404a3b25c74638d);
		test(64'h4fcf7212bebfdd89, 64'hdfd3a0870f60e072, 64'h000000002fda5ce0, 64'h5e93a0860e600042, 64'h7726ebefd8481f3f);
		test(64'h25474d793f2c7d32, 64'hb9e2a99fdb7b2948, 64'h00000004a9b27a9c, 64'h8862a8161b512040, 64'h4725794d2c3f327d);
		test(64'h0da24e08451a8d1a, 64'h44a705073f90be80, 64'h0000000003a80acc, 64'h4081040506801a00, 64'h0da24e08451a8d1a);
		test(64'h7f2e6910bdea3ffd, 64'h7fc92593c865b4c2, 64'h00000000fe552e3e, 64'h5ec90480c865b482, 64'hdf8b9640e7bacff7);
		test(64'h0f812a265e560f2b, 64'hfecee737556609f5, 64'h000000078156ebc9, 64'h4c46c226006600a5, 64'hf071da9a5191f024);
		test(64'h996d1b60923c18a6, 64'h2c1fb5204d248917, 64'h00000000026961a6, 64'h0807800048040806, 64'hd80699b61865493c);
		test(64'h4cf560811e3465c5, 64'hf2a6b292a535dc4e, 64'h000000008e485c9a, 64'h82a412100504d00a, 64'h5f3142091cb45359);
		test(64'h3b4de2fabe6d6476, 64'ha6a669d1baba633e, 64'h000000029677d59b, 64'h222660c19288032c, 64'h9d1979beaf8b71ec);
		test(64'ha73c905bcbc01878, 64'h38be984c83ce8648, 64'h0000000008f6df03, 64'h28b0000082068400, 64'h3ca75b90c0cb7818);
		test(64'h262a15662b298944, 64'hdf09e5c90a990b56, 64'h00000000068699da, 64'h4b00a0c002080810, 64'h549998a86211e868);
		test(64'ha8519a5b46242cc0, 64'h14d93f0c55095499, 64'h0000000001ad5418, 64'h0481080414014000, 64'ha765a254c01c1889);
		test(64'hbad28e0ca5854070, 64'h93d7d7a9d87056f0, 64'h0000000775314087, 64'h8142c08880001600, 64'h4070a5858e0cbad2);
		test(64'h3b0d936889b10a5d, 64'h0ec6680cabb95f09, 64'h00000000290abd2b, 64'h0206280020281701, 64'h0e3794637246ae05);
		test(64'h27429c30e8b6cff7, 64'h6465f271027abfa8, 64'h000000007126367e, 64'h64205230024abea8, 64'hb6e8f7cf4227309c);
		test(64'hd0abd7d3688aa0d7, 64'h986a686578456056, 64'h0000000006793a1f, 64'h0040482100052016, 64'hd7c707ea0ad729a2);
		test(64'hc10a152d71cb3f16, 64'h4a6c986967d5ace8, 64'h00000000849f3970, 64'h0a40980861d50460, 64'hcb71163f0ac12d15);
		test(64'h37269c228e8e3db1, 64'hf5bad73c74be6d8a, 64'h0000001e9b20677c, 64'h4120d20c40ba4c02, 64'h89cd88632b2be4c7);
		test(64'h68323fe289df33d1, 64'hcb9848f06e9659f6, 64'h00000000c4f13d74, 64'h408048b068905942, 64'hcc4762f7fc8b298c);
		test(64'h5052886f7169c8c5, 64'hb040414dd8c98a14, 64'h000000000019ecf9, 64'ha040004c40480204, 64'h88f605258c5c1796);
		test(64'hea59a91078581c00, 64'h7c6bcb08155fac38, 64'h00000000d56a9c18, 64'h3c01480000580000, 64'h001c587810a959ea);
		test(64'hbd6192029dd91d60, 64'h8a4a182923bdf75a, 64'h00000000690368d8, 64'h024818212085a600, 64'h086894e790477667);
		test(64'h8c91e2fe14041a34, 64'hc9d368e6546c1f00, 64'h00000000155df63a, 64'h8800200244041400, 64'h8c91e2fe14041a34);
		test(64'hdfd83d690e5f073e, 64'h34f2a050c605b6b0, 64'h0000000001e98f1b, 64'h20b2a000020516a0, 64'h073e0e5f3d69dfd8);
		test(64'hf3fbe985738811dd, 64'h2d21e3da342cd6be, 64'h000000013f61912e, 64'h252062100008163a, 64'h774422cd526befcf);
		test(64'h31523358d080e093, 64'hc1e3e10d162fa592, 64'h000000000a8e4067, 64'h4002000114010412, 64'hcc52c458b06c7020);
		test(64'h322721fecfeade59, 64'h4453efe0e843bda5, 64'h00000000191fbae1, 64'h0441eea060438981, 64'hfc5dde6a13b121df);
		test(64'h63c6309ca9f4f39e, 64'hb94ce939081a3df9, 64'h000000004d236666, 64'h9104e82108181c78, 64'h6df3f8566c30c993);
		test(64'h1b7769de94be57c2, 64'hb3dfbbcafb209bed, 64'h00000076eafc8af0, 64'hb1d4914ac9009b04, 64'hd7861cbabb72de69);
		test(64'h16e0c27cb6b9819a, 64'h1ab7a90d79b5d419, 64'h00000001708ccec6, 64'h08a6890860051408, 64'hbcc1d02965427679);
		test(64'hba264356875299f1, 64'h679f51136cc06082, 64'h000000000286b852, 64'h651240122cc00002, 64'hea891c592d5866f4);
		test(64'h0142aad1779780c3, 64'h3ee7342a3e84ff02, 64'h0000000004a0df01, 64'h2e66102a20006102, 64'h0418aa74dd6d203c);
		test(64'hb7e81f51b8de767c, 64'hed5fe9e149ddd590, 64'h00000015d0355f39, 64'h851c61e00998d500, 64'h1f51b7e8767cb8de);
		test(64'h1ef58a4952ff0a3b, 64'h1c4ee4e8ab011aef, 64'h000000007a85159b, 64'h1404e4e80100106b, 64'hff4adc50af789251);
		test(64'h6d8564f31f78431a, 64'ha2bd6f78450d351c, 64'h0000000051e9ce0e, 64'h00bc6c10000c0508, 64'h3f4658d6a13487f1);
		test(64'h896063c58085e876, 64'h40f7cd92ebbc3e26, 64'h00000001826411a7, 64'h40600400ab201c24, 64'h02522b9d6209c953);
		test(64'h8fbe5684b9140fda, 64'h7daef51856149145, 64'h000000000ff584cc, 64'h3882400056141104, 64'hf4d79a846782f05e);
		test(64'h6a01074de3fa4927, 64'h9ef4f552e7611475, 64'h00000001401cef0b, 64'h8e84f51042200415, 64'h68b13d5fb0e85920);
		test(64'h298564256e5e6b1d, 64'h10f1368a1f6db08b, 64'h0000000011a0eb25, 64'h1070128a064c1089, 64'h1a494a62a7678b6d);
		test(64'h5d56f9d1347a292a, 64'h8ea99d9b624dd7f8, 64'h000000060ee56025, 64'h0209109a40091150, 64'h2a297a34d1f9565d);
		test(64'h34023e3619adb257, 64'h9ad02588915e9cf3, 64'h0000000010619b17, 64'h1850048811188453, 64'hd4ae895bc7c6c204);
		test(64'h74c5fd46fe517d0a, 64'h3b68686e72b3dd70, 64'h0000000313cfcaf8, 64'h2b68404822b28120, 64'h7d0afe51fd4674c5);
		test(64'hece19f6bb49be6ca, 64'h3ee4838f7edc2387, 64'h00000005bbadab6a, 64'h1cc401067c542082, 64'h3787f9d62dd96753);
		test(64'h22d0e03f67599a00, 64'h7b315baeaed9a934, 64'h00000004941eb7d0, 64'h79205928a2900000, 64'ha90076950ef3220d);
		test(64'h5e36e6f8de04d766, 64'hde684601baf1c748, 64'h000000001f5d707e, 64'h5c0002003270c140, 64'h365ef8e604de66d7);
		test(64'h947f5b84d090f6c6, 64'hc3da19bcae82a6ab, 64'h000000010ff185f2, 64'h42801080ac82240a, 64'h90b036f6ef9212ad);
		test(64'h2f041032f1ef6926, 64'h397e4f777e1a3e74, 64'h00000058406b8745, 64'h182e41736c102430, 64'h96621ffe0123f240);
		test(64'hf29b22bb7fb71708, 64'h3c4fd90e7020bb26, 64'h000000003160be58, 64'h3c4d990050208100, 64'hfdded4208fe688ee);
		test(64'h50a82c31942af3d0, 64'hd097050107aa5237, 64'h0000000001c2c7e8, 64'h00120401070a5020, 64'hcf0b2954348c0a15);
		test(64'ha728015173d16b53, 64'hf0a63b79f28c7d45, 64'h00000005206af9ad, 64'h20a41b20b0845405, 64'hb541202a3b2e793a);
		test(64'h19e2cc9f042094ff, 64'hdc778f6734be0a16, 64'h00000001b2e1ca07, 64'hd0040402108e0a16, 64'h33f6648b16ff1008);
		test(64'h9386770d73133382, 64'h7066804ea183b565, 64'h00000000013336d0, 64'h3002000c2101a004, 64'h3b3233143694bbe0);
		test(64'hb483dfd4bc1f4b4f, 64'hbb684d7f77ee4619, 64'h000000381f51c1eb, 64'h28484c0764aa0219, 64'he8ef43788f872f7c);
		test(64'hea295863c3f93cd5, 64'h141ed10a6a735bec, 64'h0000000008ccf599, 64'h1002d10a08330aa4, 64'h9f3c5dc392ae3685);
		test(64'h095af16505bac65b, 64'h2d3b4ee773e54517, 64'h00000005743a1a6b, 64'h0900466530604113, 64'h8fa6905a63daa05d);
		test(64'h9bdbb638b84b2a5d, 64'hdc21e506a8288b49, 64'h0000000002cd8eb7, 64'h0801600488008341, 64'he76734798774ae15);
		test(64'h85874e05ee0d281f, 64'h94d8fb126886d58f, 64'h00000000b098e80f, 64'h945803020804008f, 64'he1a1a072b077f814);
		test(64'h0c70adc8009b5be4, 64'h64fb84e0f5961453, 64'h00000000171e0368, 64'h0008846054961010, 64'h5b3103e0ad72009d);
		test(64'hbe8273820a044cbb, 64'h5c5ddb8f13500ae2, 64'h00000000381b922b, 64'h0410080910400aa2, 64'h0a0113eeeb28dc28);
		test(64'h25cfd1c67cc65277, 64'h3e8ce7a94dc3a313, 64'h000000012f8c7717, 64'h0e8860a04440a213, 64'hb8364a3fa4eee336);
		test(64'hd8270a281af88095, 64'ha3db049a0d57f4d4, 64'h0000000080c5310b, 64'h0193049004004444, 64'ha0828d720859a18f);
		test(64'h69bbf1ef4e50ee3d, 64'h3f832675d87260a1, 64'h0000000029f36b5b, 64'h0e02201558026081, 64'h8da0dd3e9677f2df);
		test(64'h5779c0dc7b0e8c20, 64'h79f9289de3af9938, 64'h0000000abe79e754, 64'h60f12005a0281000, 64'h208c0e7bdcc07957);
		test(64'hdfd0c092d0bd880a, 64'hf92dc94f084bb19a, 64'h00000000dc304583, 64'hd004c90c00400088, 64'h6830707f0a22e770);
		test(64'h00a9c51ef2760079, 64'h26b72b5d366fd239, 64'h0000000188bb760f, 64'h2636085920005221, 64'hb600b9f12dca5600);
		test(64'hab4cefeaaa0aa3dd, 64'h85618ac56a39e1da, 64'h000000002cf8e57e, 64'h812000412201e0d2, 64'hbabf13ae77ac0aaa);
		test(64'h1ecbf0901b9ca499, 64'he010d0277f319b90, 64'h0000000000e06d43, 64'ha010802629010a10, 64'hf0901ecba4991b9c);
		test(64'hd49d8a08f7951ca7, 64'h3eb06c805e15ff5e, 64'h00000001549be383, 64'h0e9068004a00e50e, 64'h20a27617da3456df);
		test(64'h7c5eeff7e27dc320, 64'h07dd06c4cbe1f0a6, 64'h0000000047bfa7c4, 64'h061106c0c8212000, 64'h8b7dc3083db5fbdf);
		test(64'h8f449cba3190dac7, 64'he69008066ff9aab2, 64'h00000000265464b9, 64'hc09000020368a032, 64'h7a3dc46063ea2f11);
		test(64'h2ebab447c2d4b567, 64'h29c8f524254aa5cd, 64'h000000001adc89eb, 64'h0088a4040508850d, 64'h57d1b8878e1cb9a7);
		test(64'h65de7f4fac9ce3c6, 64'h60f0f4c25f87eb81, 64'h00000000f5ecccee, 64'h40b020c20e03c180, 64'h9aedbf8f5c6cd3c9);
		test(64'ha20de1288f9e2416, 64'h5c615a2f4636ddde, 64'h0000000018c3708b, 64'h04005a234404404c, 64'h284b708a9418b6f2);
		test(64'h80d266e0417c07e5, 64'h29b2ce151357a6aa, 64'h000000000b583c3c, 64'h20024e100007a422, 64'hd314b50d7820b099);
		test(64'h69debc3cde83e367, 64'h946362f6c168dd61, 64'h000000000a47618f, 64'h84624016c0089861, 64'hed43d39b96ed7c3c);
		test(64'h7a911b4c8447749b, 64'hacecbed09b65bcb2, 64'h0000000681aa16db, 64'ha080841093442492, 64'hd16e211d4e13da64);
		test(64'hba8e69b3623c1b4b, 64'h9ca964d0abedd1bd, 64'h0000000756aa38c5, 64'h18a02010a80cc115, 64'h7872c3193769d457);
		test(64'h9fcf80bdc145c55e, 64'h7ecf2edfe1b5d954, 64'h0000003ff0bba3cf, 64'h5e4c0242e0114950, 64'h08dbf9fc5ce51c54);
		test(64'h6cbbeb1847e667e6, 64'hb5bdd63a675e92a9, 64'h0000000af72d799c, 64'ha021d60a061e9028, 64'hd98bd99b779c24d7);
		test(64'hd0ac43275df9a5cc, 64'h2beb8aec129ca587, 64'h000000000b096efc, 64'h09cb8a281014a084, 64'h0b35c2e4ba9fa533);
		test(64'h935e96eec3381d0c, 64'hd129ee258f74ae36, 64'h00000002d47a6c62, 64'h9100622400708030, 64'h7430c32c96bbc6b5);
		test(64'he7dd9c7a99530aea, 64'h8166d932f500567f, 64'h00000000756f28ea, 64'h006091028100126a, 64'h5750ca995e39bbe7);
		test(64'h57cfb2fd88162913, 64'he72244a4f0ac2181, 64'h0000000000ba781d, 64'h0222002090040081, 64'habcf71fe44291623);
		test(64'hc0e19bee65713982, 64'h2da6ea653427fb71, 64'h0000000064fac9d0, 64'h28a0a26010073010, 64'h36419ab267ddc0d2);
		test(64'hc1fb89c6995148c7, 64'h09100e0b1e053b96, 64'h000000000071624b, 64'h0100080212001816, 64'h629343ef21d36645);
		test(64'h96e0931a06c71461, 64'h2d4017622591a209, 64'h000000000016caa1, 64'h2040142020110001, 64'hd0692563cb099228);
		test(64'h391c6891f7e9230d, 64'h20e65e9f2e39920b, 64'h00000000454c6ecd, 64'h20c65c8420300209, 64'h83c9986179fe0b4c);
		test(64'h4abe88aeab9e03ef, 64'h8c51a90e99642428, 64'h00000000004abd93, 64'h8051800019602428, 64'h9eabef03be4aae88);
		test(64'h8dae2963951ae660, 64'hf6fdcffddf1d4bac, 64'h00001156258d5ca4, 64'h44c585454e0c0a00, 64'ha159066eead83692);
		test(64'hae70e5fe7ef21a3b, 64'hdb424fe85c5010cf, 64'h0000000026abffcb, 64'hda424900540000cb, 64'h0e757fa74f7edc58);
		test(64'he64f0f005ca9632e, 64'hb298eec62efd3a68, 64'h0000000691c1aacb, 64'h0088c4840a8c1260, 64'ha95c2e634fe6000f);
		test(64'hf881de090e9b5a1c, 64'h3e8ddc0306436ba8, 64'h000000001c9fbbb1, 64'h1c81980206020380, 64'h9b0e1c5a81f809de);
		test(64'hcb625c72f31e077f, 64'h35c7f93918f404b1, 64'h000000000a96c877, 64'h3444780008d404b1, 64'h0bbff32dacb1c791);
		test(64'hfc52b53616a2e0f8, 64'h95ba835cb85a9b39, 64'h00000001c5aa430e, 64'h0098810438001b20, 64'hf4d05129397aa1fc);
		test(64'ha8a43fa8c475c04f, 64'h25dfe461809ad80f, 64'h00000000244354cf, 64'h008744600000400f, 64'h251515fcae23f203);
		test(64'h3f550f8222d20e7f, 64'h9d07a6f8789dd5a3, 64'h00000003e9c13027, 64'h100422a0400d15a3, 64'h44b407efcfaa0f14);
		test(64'h587b33e3d83de6c8, 64'hb2901e2ff2272f05, 64'h000000001333d6d8, 64'h9200022de0252200, 64'h4a7b333d4ee39d4c);
		test(64'h2760c87bc1de001b, 64'he0526c9d3468dadb, 64'h00000000329a280f, 64'hc0002c1d00000053, 64'hed31604e8d00b738);
		test(64'h3f92575fb431ddae, 64'hd0a72bac17b11595, 64'h000000001919e3fa, 64'h50200a0c13910494, 64'hbafaf316eed58723);
		test(64'h2da80edbe495b2fe, 64'h057014720c59e61b, 64'h00000000034dab5e, 64'h004010520441661a, 64'hbd07514bf7d49a72);
		test(64'h55542ca5a4d5b317, 64'he37fc02b17f03db1, 64'h000000026a129b93, 64'ha249802215902131, 64'h732b58ea1c5aaaa8);
		test(64'hb46d235d9972918a, 64'h2a80c4f980875629, 64'h0000000001017922, 64'h228080a100030208, 64'hb16645629e78ae13);
		test(64'ha47aba2d5d1cf2c5, 64'h2d82d2286a02da60, 64'h0000000000a6fa76, 64'h0182122808028220, 64'h5d1cf2c5a47aba2d);
		test(64'hd685928e6e8447d4, 64'h8bdd40842f043a5b, 64'h000000000a8dfa38, 64'h8a81000021043848, 64'h17941ab6b22e1267);
		test(64'h9e569cd1e8c1c4ef, 64'h3c43bf737ab09ca6, 64'h00000003eb95d49f, 64'h0c428601608098a6, 64'h2b4313fbb6953647);
		test(64'h5c30cc690bc8141f, 64'h68a2c478eeb763f7, 64'h0000000abe8b000f, 64'h4080043888024037, 64'h28f8d01333963a0c);
		test(64'h34773f857f2c10f0, 64'heca0e6d0d56a74d1, 64'h000000002a78f62e, 64'h6ca084c001007400, 64'h3f4a38bb20f0bf1c);
		test(64'he290c80a0837b478, 64'hae5b64956d65c510, 64'h00000000651008f5, 64'h040144946405c000, 64'hc80ae290b4780837);
		test(64'h761b167333584a9a, 64'ha10cce0633611c8f, 64'h000000000286fc5a, 64'h210448002120108a, 64'hd86ece681acc5952);
		test(64'h184819d8fe3d1d76, 64'hdb63264296b0facc, 64'h000000003205ec65, 64'hdb40264080b05a48, 64'h84818d91d3ef67d1);
		test(64'hfa2f6388f088a839, 64'h94b76debf8169729, 64'h0000000cbe64f087, 64'h80360420a8000701, 64'h44f036541ff54493);
		test(64'h7461f78058285047, 64'hf4fc6e75bacaf127, 64'h0000003d8d80c4a7, 64'h0014402408802007, 64'h1a140ae22e86ef01);
		test(64'h00fdc6d1272dcd05, 64'he2b64290180e77df, 64'h0000000007bcd285, 64'h40b04090080c3205, 64'h8b63bf00a0b3b4e4);
		test(64'h389463a20cb87cf0, 64'h716b303109323009, 64'h000000000030296c, 64'h3101303001320000, 64'h68345193740cf0bc);
		test(64'h8129086f8dff7629, 64'hc12337db86f62285, 64'h000000005a05f7f9, 64'h002237d984c20201, 64'h246140f9e4ff9b61);
		test(64'h498167ccd723cf80, 64'h7c17f3ce2fb0681f, 64'h000000090b7e3aa0, 64'h6412e10629b04000, 64'h33e6819201f3c4eb);
		test(64'h57c24fb98ce8ef0f, 64'h37b8a48ee2091d11, 64'h0000000007c1c89d, 64'h31a8008ce2000511, 64'h8f76abc1df0f4cd4);
		test(64'h7713966e88fe6b6b, 64'hf22ab5cffde22d7d, 64'h00000079b3d13f75, 64'h62288107f1a02955, 64'h7979df44d99632bb);
		test(64'h7c14d29d73f31667, 64'h03be5c21c40b898b, 64'h0000000000562983, 64'h01bc18008408880b, 64'h82e39bb4fcec6e86);
		test(64'he979f8c8cce09c58, 64'h96e0cd3ce0154b60, 64'h00000000087c2c12, 64'h90e00024c0010a00, 64'hcce09c58e979f8c8);
		test(64'h3161b44b4607b9f6, 64'h1d824184b0510b05, 64'h0000000000120036, 64'h0582018410510904, 64'h2329877898b0679f);
		test(64'h315aaa061cb5c853, 64'hde5554aa2af2d703, 64'h00000000460156c3, 64'h0641142228404403, 64'hc8a5550683da31ac);
		test(64'h5786a032bc28926d, 64'h6e36742b312bf809, 64'h000000004cd2b64b, 64'h2e0050021008d801, 64'h49ab3150147c9e61);
		test(64'h49a6d14749c48db9, 64'hdab76b89b2074ae2, 64'h00000000ada2422a, 64'h9087020812030a82, 64'h163127e616a9741d);
		test(64'h954c42a9b003bcf7, 64'h91a26e64588e664e, 64'h000000001c45216b, 64'h800000641888660e, 64'h31566a81c00edf3e);
		test(64'haca8c6612d6b2902, 64'he11b8bbc2f7bffd0, 64'h00000052523bb948, 64'hc002099425492040, 64'hc661aca829022d6b);
		test(64'h3dd33a0e0e7efc2f, 64'he64b7a878676ea17, 64'h00000001adecffe7, 64'hc0034a8706740817, 64'h5c70bccb3ff4707e);
		test(64'hf2b22e590d846203, 64'h4dfb587946c98a07, 64'h000000008b46ea0b, 64'h00d8080900800003, 64'h4f4d749ab02146c0);
		test(64'h163bf68dc6c078d3, 64'h5da95e5a3b8dace2, 64'h000000029f64286d, 64'h4d014c000b80a422, 64'h3930d27c49cef927);
		test(64'hccbd6f02477bcf3b, 64'h5ada5461c82b9665, 64'h000000002ad42fb5, 64'h02ca5061802b0645, 64'hb87bfc73cce7f910);
		test(64'h930a269b8380f809, 64'h1efa7337fccadbb9, 64'h00000121a9704783, 64'h08da003404ca0021, 64'h06f4404367190563);
		test(64'h3b524052fa6e804e, 64'h2dfc874609af8ece, 64'h00000003540b3d0f, 64'h25e806460100044c, 64'h85ec8501b9afb102);
		test(64'h619051f25b20a253, 64'he63f814b4c5a17d7, 64'h000000018835809b, 64'h8436010008401143, 64'h8a4f860945cada04);
		test(64'h9c19d86ae2cdb638, 64'hfc2cc87e740aa354, 64'h000000004ebeb972, 64'hc40c085a54002300, 64'h8da6c9916b832edc);
		test(64'he40cfcb31804e312, 64'h2e746c503fc66e54, 64'h00000000a1f582ca, 64'h024000100e060410, 64'hcf3b4ec03e218140);
		test(64'h8c46d0ae4cf8f788, 64'h28f9de58f863e467, 64'h00000002870539e0, 64'h28218e503843c020, 64'h321fef1131620b75);
		test(64'h5ab8ff1b9938da6f, 64'h3398cdc75b47d01b, 64'h00000000dfe36877, 64'h309041c05304c01b, 64'h8dffd1a56fb5c199);
		test(64'he7b19aee8cf0397b, 64'hf2894677a55ae7c9, 64'h0000000769dab097, 64'hd001407400584789, 64'h72dbdd65f04cb736);
		test(64'ha081bd1840dc8046, 64'h76df5e8206f9e8c6, 64'h0000000220b83687, 64'h02014e0004004044, 64'h0a427e2401370291);
		test(64'h9cf6034c54b8ea97, 64'h31b7483b427dde82, 64'h000000005f049cd7, 64'h1091083042548a82, 64'h63f90c1351e2ba6d);
		test(64'h596960899b20c5bf, 64'h3306126a4f780bf4, 64'h000000000a04b437, 64'h310402000c2809f4, 64'h5cfbb90206989596);
		test(64'h6acd4407495c86e3, 64'haf2436114e6fe72e, 64'h00000001a49cb269, 64'ha42012014841a606, 64'h3561cb9273a9d011);
		test(64'h8e73c43d6d2f3360, 64'hf58ef5e0d059b506, 64'h0000000110e451b4, 64'hb1845580c018a000, 64'hb2cd137c79f8cc09);
		test(64'h3f0ce85d3eec87ec, 64'h217c1f85e48b25e3, 64'h0000000063433c7c, 64'h01781d80800b2560, 64'hc7731e73cf0371ab);
		test(64'hd76ce83cffe72b68, 64'h08a09451e4c33f3e, 64'h000000000317fd74, 64'h08a09440e0411b10, 64'h29e8dbff3c2b39d7);
		test(64'he12edddd7da2b6c0, 64'h8bfbaad57e7643ad, 64'h000000496affc950, 64'h83aba2902a544200, 64'h15eb0c97d12deeee);
		test(64'h717f45ce49bbe46a, 64'h9b348f595518c922, 64'h0000000009e5a9f3, 64'h11248b5810088820, 64'h16eeb19ad4df153b);
		test(64'h3fa96bf858c4f030, 64'h8ab1c2bfecef75d0, 64'h0000000f5f8564e1, 64'h8801420c44e01400, 64'h6bf83fa9f03058c4);
		test(64'h553b7ffff827df3b, 64'h2944e274894d3e45, 64'h00000000023fe379, 64'h20004074814d0e05, 64'haa73fbff4fb1fe73);
		test(64'h7b174e0abe2a9579, 64'hf80b53450f7abe13, 64'h00000000f7439755, 64'h580b01040a289e01, 64'h2705ed8e9ae9d745);
		test(64'hf9d92d5c5357afaf, 64'h593bd5a6dd8f0b30, 64'h00000003da3264fe, 64'h01119126958d0330, 64'hafaf53572d5cf9d9);
		test(64'h03de352aa0dcd926, 64'heb1724ec8ba7e914, 64'h000000001f668a6d, 64'h480120e089824110, 64'h53a230ed9d620acd);
		test(64'h4e732c2381e463c6, 64'h4eeed5a806859a81, 64'h000000001ec89186, 64'h00e8818002850280, 64'h8db31c1342d893c9);
		test(64'h50d7ebae675611f4, 64'h6aed3b4ead8c40d7, 64'h0000000233bbacbc, 64'h428d1248080c40c4, 64'hd7750aeb882fe66a);
		test(64'h025a5099c0f18d96, 64'hbc74071568bbcb0d, 64'h00000000050b39aa, 64'ha00407006019820c, 64'h5a10660a2f0c96e4);
		test(64'h3243aca5aa4fdfdb, 64'h28e7a5f0245fd6a4, 64'h0000000093eaaffc, 64'h20a220f0241fc624, 64'haaf4fdbd2334ca5a);
		test(64'hf9934055a9244009, 64'h1d8d405596f52ac9, 64'h00000000367f0503, 64'h1408400404000081, 64'h63f6aa8018560680);
		test(64'h4e30b6f8807352dc, 64'hab287642010e8379, 64'h0000000000d3e156, 64'h0320320200048270, 64'heca1b340f479308d);
		test(64'h48b5db89d6bd603f, 64'h231ae4032c31f53f, 64'h0000000004c4f63f, 64'h0218a4030830003f, 64'hfc06bd6b91dbad12);
		test(64'h166985e06a993915, 64'h61dc75e3f76eee27, 64'h0000000a1f1910c5, 64'h61003142622c4205, 64'h56999ca86896a107);
		test(64'h788ea6e682895a3b, 64'h09bf5f618a03a64f, 64'h00000000a70daa2b, 64'h080504410a01024b, 64'h711e67659141dc5a);
		test(64'h726cb29218b1d2c3, 64'hfd38d93fe9e061a6, 64'h0000000716890ac9, 64'h20301123a0a04006, 64'h244e87c38d398e86);
		test(64'hd344de75f3d508e5, 64'ha185ec173b043bb4, 64'h000000002adeee4d, 64'ha005c81202001a24, 64'h805e3f5ded573d44);
		test(64'h16fda375ee8c5ec3, 64'hd2e463a400e296be, 64'h0000000007eee1e1, 64'h5240220400628606, 64'hc3b532bb5dca7f94);
		test(64'hdad3875d5ab73c13, 64'h13cb08cdc71936ab, 64'h000000006d9eabc3, 64'h118900c583180083, 64'hdea58cc3bcb5ab1e);
		test(64'h58aa6d512003ce06, 64'h86adbf22eb44881a, 64'h0000000007168419, 64'h8000072068000018, 64'h5497aa52093b0c80);
		test(64'hd236ace861a7478a, 64'he89e9714674eab85, 64'h000000018ba1931c, 64'h28028414440e8104, 64'h1e93c54d29b5b854);
		test(64'hfd9c717ea67e7792, 64'hf6a0d64055a72ffd, 64'h00000007d324ebc8, 64'hd200c24055070f24, 64'h16bbdb95db2bc6ef);
		test(64'hf72abf3d24fc3ee2, 64'ha2a74d599a583e1f, 64'h00000001d4ee1fe2, 64'h80820d5802582e02, 64'hbcfd54ef477c3f24);
		test(64'h864717af6be6e9a3, 64'h5a37bc5848df2cb0, 64'h000000001394f9b6, 64'h1827a44848462030, 64'he9a36be617af8647);
		test(64'h34b5980e57c1bee9, 64'hf21c23eac374a7d4, 64'h000000006a06f1ec, 64'h220c2300c1742684, 64'h89e0435beb9e751c);
		test(64'h046b073128173b9b, 64'h14ab69828ea2932c, 64'h0000000002f110ba, 64'h000129008ca2030c, 64'h7182b9b3b6401370);
		test(64'h6524ecdb4b6a9d0a, 64'h0c341349e19a4ab0, 64'h0000000000d1d4d0, 64'h0830110861100220, 64'h9d0a4b6aecdb6524);
		test(64'ha5092e1ff9d7d225, 64'h08c5d7afe01654c1, 64'h000000000118fff1, 64'h0881c5ad20004081, 64'h5a061d2ff6ebe11a);
		test(64'h24a0aa4ca08b6828, 64'he9c8000b9fe574f8, 64'h0000000012482385, 64'h400800008da00440, 64'h28688ba04caaa024);
		test(64'h2a3b5f21df3a8011, 64'hf542de42a084d151, 64'h00000000010be443, 64'he142480000001001, 64'haf1215374022ef35);
		test(64'h915aa2f1c7bdacb3, 64'he2ea6ead489b9b2a, 64'h00000002169cdda5, 64'h620a66a508188a0a, 64'he73deca35a64f4a8);
		test(64'hde0337230ab1269c, 64'h882510a5039c63d1, 64'h0000000000cd6c6a, 64'h80240020021841c0, 64'h3b13ed03196c0572);
		test(64'h8d0b96443c558f56, 64'hd1e6b6a5733431c8, 64'h0000000090dc98ca, 64'h11c09224132410c0, 64'h0b8d4496553c568f);
		test(64'hfed8993c25b12bab, 64'h2b46ca3a92bdc33c, 64'h00000000e95c393a, 64'h0204c2208095822c, 64'hbab21b52c3998def);
		test(64'hc55e7a421ffbf7ba, 64'h219e22534664aed5, 64'h000000000bfa7b74, 64'h219e22434644aac4, 64'h5b18acdabf57f27f);
		test(64'h200a3a38098972c8, 64'h257dca4091c5d22d, 64'h0000000010431974, 64'h043082009104c020, 64'h64604c1b50014353);
		test(64'hfa9c04663e4572c9, 64'hbeb7785119e46a6c, 64'h00000003db0265da, 64'h86b1081019206044, 64'h54e39c27c9af6640);
		test(64'h12a8beda3cf0b9b8, 64'h38145996ce0636cb, 64'h00000000086d3194, 64'h380059008e0032c0, 64'h5184b5d7f0c3d1d9);
		test(64'h28ed84cb7402e866, 64'h9e7b7d27d7303436, 64'h000000026a11b84b, 64'h8c720005c4003014, 64'h2b991d8012e3287b);
		test(64'h81a09ce561a999de, 64'h027bacdf08ed7d6d, 64'h00000002179569b6, 64'h005300ca00c51c6c, 64'h6529de660524adc6);
		test(64'h6dbdc9459ba05cd7, 64'h74b7b6f06046c9ae, 64'h00000001bec100d3, 64'h60a720102044488e, 64'h0ae6d7357e795163);
		test(64'h5077f98e977befbd, 64'he076f585871d5722, 64'h000000005ff77ede, 64'h80567485851d1702, 64'h6ddebfe750ddf62b);
		test(64'had620aa92bbae50c, 64'h6eecd66b6c7953c6, 64'h0000000e605ace92, 64'h222454692c1100c0, 64'h7a89a06ae8ae5b30);
		test(64'h04eee588af4f90e1, 64'h46ec7053b0e91780, 64'h0000000005fc1971, 64'h46a0705080290080, 64'h04eee588af4f90e1);
		test(64'h5df3d438446325af, 64'h4d20a42398df6824, 64'h0000000003f6046b, 64'h01200022104d2824, 64'h443652fad53f4d83);
		test(64'h643b94f6bad85ff4, 64'h04dddda3ced2924b, 64'h0000000136aeaf38, 64'h009c998046d29208, 64'hcd62f692b1d5f2af);
		test(64'h5075a874e4fcc5af, 64'h61b497e1c579b7e4, 64'h0000000478377a5b, 64'h40b011e1814132e4, 64'h4ecf5cfa05578a47);
		test(64'h8e8ee2d415743d8b, 64'hc305077bc980d730, 64'h000000000a950234, 64'h41010641c8808230, 64'h3d8b1574e2d48e8e);
		test(64'h3643233771fc1a9e, 64'h5fa44007e91c852b, 64'h000000000583b786, 64'h07a440002814012a, 64'hf3e897852cc6ce4c);
		test(64'h3eb796cb1c8896e1, 64'h9c975c2085501f8c, 64'h0000000003fd48b4, 64'h8402080081401c04, 64'h7be3bc6988c11e69);
		test(64'ha3da4d4a2acadcb3, 64'h37a1417f5c2a05ca, 64'h00000000273944e9, 64'h252100565808050a, 64'h7aac1a173a8aec73);
		test(64'h70ee66fb2e286341, 64'h7f39dd31d98ac3c7, 64'h0000001c292e24e9, 64'h6c29842018028201, 64'h0e7766df7414c682);
		test(64'hf78fd82f0ff1c780, 64'h57d6077d1d71c40f, 64'h00000003f30bbff0, 64'h5056074510710000, 64'hf1eff41b8ff001e3);
		test(64'h3922d0ed0b35c447, 64'h7d2846dc18c45e0f, 64'h000000001da6d327, 64'h1500449c00400807, 64'h449cb70bacd0e223);
		test(64'h3186160870c5b573, 64'hdee059eee25502d9, 64'h0000000044411acd, 64'h1c00504cc2110289, 64'h04294932b37acab0);
		test(64'ha9282bbb77b23e9c, 64'h5a88afc551c37de1, 64'h000000004b73e9e8, 64'h4a80ad8100c351c0, 64'hbb713d6c56141777);
		test(64'h84036df182b7a35a, 64'ha656577e8d095a9c, 64'h00000001435e2116, 64'ha002133c80091288, 64'h1fd63048a53a7b28);
		test(64'h87c4c7fec7446f29, 64'hcd55a5407d5a0db7, 64'h000000013abc71d1, 64'h48152000451a0891, 64'hf694e322e37fe123);
		test(64'hda738494824d346c, 64'h065debe6f4813504, 64'h000000001cc1283d, 64'h00088a8640811400, 64'had37484928d443c6);
		test(64'h546f0817d359f66e, 64'he7370106284b1e02, 64'h0000000000a5d9b7, 64'ha307010428030e00, 64'h519f024d7c56f99b);
		test(64'hd01741bfc46048be, 64'hc8d3ad9b65b367af, 64'h00000031c3fa443e, 64'hc8d3040a002102ae, 64'h06237d12e80bfd82);
		test(64'hbd44a60746140aa0, 64'ha567dfc559a48ab5, 64'h00000007d231c178, 64'ha441828001208200, 64'h5005988295b0e788);
		test(64'hca121cdfb6a3cee0, 64'h7b25481dba1b317d, 64'h00000001307fa630, 64'h6a244010b80b1140, 64'h0ddc3597fec2125c);
		test(64'hb6c271b99132f85f, 64'hab354a52257b6a6f, 64'h0000000341116baf, 64'h28204050047a022f, 64'h4c89fa1f436d9d8e);
		test(64'he3ba95ad7c50e77b, 64'hf8cb78aede94f875, 64'h0000003962f3cb9d, 64'hb08b60240e04d865, 64'hbd7bcb0aa6e53d57);
		test(64'haa846c0860936cc5, 64'hf2ff18f98fa9db5c, 64'h000000ac22102549, 64'h020c00480d891814, 64'h80c648aa5cc63906);
		test(64'hc37eb209127fdfea, 64'hcbd927c551fb9ad5, 64'h0000001b750a7ff8, 64'h410804c551db9a44, 64'h17603cdbfe5d12fb);
		test(64'h733c632927a478a0, 64'h1403d29023431851, 64'h000000000010a718, 64'h0002129000410000, 64'h9316b33cb4501b58);
		test(64'h842614c6e48baa21, 64'h2dbdc81f14861535, 64'h0000000009206689, 64'h2110881a10800401, 64'h55218d74829c8491);
		test(64'h3822c5c32132f45f, 64'h4916fe2a79a86677, 64'h000000011c452baf, 64'h4804122059880237, 64'h2ffa844ca3c31c44);
		test(64'hbb048165dd7a4b7b, 64'hfe0068c50367012d, 64'h0000000002e8775d, 64'h5e00204002630125, 64'h5bee7b788077a924);
		test(64'h008f9830f85a246f, 64'hda0503691c606be7, 64'h0000000000c4d21f, 64'hc0010148040041a7, 64'h1f5a24f600f1190c);
		test(64'h9bd546d9bedeb2f0, 64'he8a8b5430b7bb395, 64'h0000000130575dec, 64'hc8a8944309313300, 64'h986e76ae170fd7de);
		test(64'h54f49e62269701b2, 64'h90bde55da14e0331, 64'h000000001ea5046e, 64'h80344540004a0210, 64'h0271196b6d91a8f8);
		test(64'hd7e36e026f047377, 64'h701d2cf5a80a4651, 64'h00000000051e032f, 64'h7000083428024451, 64'h9d01ebd3b3bb9f08);
		test(64'he9a68cc4c43be69d, 64'he898175813b99610, 64'h0000000007c481f7, 64'h8018135801909410, 64'h8cc4e9a6e69dc43b);
		test(64'h0dad0d77bd41613c, 64'h570fa1a277b82cfe, 64'h0000000174b7421e, 64'h560f208005800878, 64'h3c49417edd707a70);
		test(64'h936a290c9e8da327, 64'h8cb60cd1b3fe91a1, 64'h000000008982d1ab, 64'h80b40811311880a1, 64'h6d4e531b6395160c);
		test(64'h880018c9748d24c2, 64'h8267c75efda34e0b, 64'h000000040051d492, 64'h0047410648814002, 64'h001139811be23442);
		test(64'h7bcf824e95e4ea57, 64'h3236852d40395643, 64'h00000000039c644f, 64'h1230802c40104443, 64'hed3f14279a7275ae);
		test(64'hf5b67739967ad42f, 64'hf5dda5b0b5e8ca47, 64'h0000000fea7767c7, 64'h944c259031400847, 64'haf6dee9c695e2bf4);
		test(64'h893e0b9963df6a13, 64'h33872aad2b8e3007, 64'h0000000002ceb7f3, 64'h01862aa509002003, 64'h917cd099c6fb56c8);
		test(64'h82f98268cf1bcda7, 64'h56a8b138463a73fc, 64'h000000001f17bc69, 64'h50a880304622529c, 64'h7adcb1fc86289f28);
		test(64'h0d174a260663781b, 64'hbe64569a0de4d82b, 64'h0000000018c8a677, 64'h024050180d800823, 64'h6c068de18e0b4625);
		test(64'hc6cfce902d7a7b5b, 64'hde31c9036e0f396d, 64'h0000000199e1d5f5, 64'h0a214902460d2865, 64'h5be17a7bfc9c06dc);
		test(64'he9c99feab48edc5f, 64'h9a53935ff5953627, 64'h0000000a9faaea67, 64'h88431043b1901227, 64'h2d713bfa9793f957);
		test(64'hd3850ed862e1758b, 64'h0fb837102f88b5a0, 64'h000000000383653e, 64'h02b002102a8804a0, 64'h62e1758bd3850ed8);
		test(64'h0441701962d8cccb, 64'h9be32794a0932f92, 64'h0000000001309c65, 64'h90a2241400902912, 64'hd0460114333e9872);
		test(64'hdf2c01369271ad4d, 64'hd2086bf12c39bd57, 64'h00000001f0986ef5, 64'h400808e00c119415, 64'h806cfb34b5b2498e);
		test(64'h9b1d4da2007e7bed, 64'h8da1768d2c29dc5a, 64'h0000000069940cea, 64'h000036882c21d852, 64'ha817476eb7dedb00);
		test(64'hc76a3db5b549d962, 64'he5c85cf813d95250, 64'h0000000036ded57a, 64'hc488087012490040, 64'h3db5c76ad962b549);
		test(64'h0ff78ffed60874f4, 64'h74df0bda151dd91d, 64'h00000000f7ffc8ca, 64'h6496004005145908, 64'hdff4bff08f8b409e);
		test(64'h9759bb2f56bc05ef, 64'hf3ca6600ebe5e624, 64'h000000009d952b0b, 64'h518866000045c624, 64'h65cb50fe7995bbf2);
		test(64'h61613094e65f24e8, 64'hd1f23288fd85a0a1, 64'h000000000acd726e, 64'h1122328048852000, 64'hd9af18d492923068);
		test(64'h404819677e42a3a0, 64'h3d66d787e9accee7, 64'h0000000209770468, 64'h3162d60421204c80, 64'h7e42c505021298e6);
		test(64'heb972fc689e4ceba, 64'h4c7ce920375de9a7, 64'h0000000314e0cb5a, 64'h440869001145a1a2, 64'h9127735dd7e9f463);
		test(64'h6cd264efaa15dbb4, 64'h3d13980d71479d03, 64'h0000000016c3a2f4, 64'h1400880551071900, 64'h63b4627f558abdd2);
		test(64'h6a1d818dac1032f9, 64'h03570650aca38cdc, 64'h0000000004d0f01e, 64'h020100000c028cc4, 64'hd818d1a69f2301ca);
		test(64'hb19c80e7ad087cc5, 64'hca9b2a07d52dfd7c, 64'h00000008e0f347d1, 64'h4a892200400dcc14, 64'h5cc780da7e08c91b);
		test(64'h60823baddd5b7986, 64'hf9b5111862e56ef5, 64'h00000001886c4f22, 64'h71a4101822650c14, 64'h6b94ee7a73e50914);
		test(64'h39ddbc353475b968, 64'hd65a4432e46a081a, 64'h00000000009ce3ca, 64'h0648441284280800, 64'hc5e377c692e6d5c1);
		test(64'hdefc14c9ef379a8a, 64'h9a2767c16c20173f, 64'h000000007e13fe8a, 64'h922625c10c00120a, 64'h5159ecf793283f7b);
		test(64'h9f913ce515b878d1, 64'hb3a0f84086571c60, 64'h0000000002f1e91a, 64'h31a0084084061020, 64'h15b878d19f913ce5);
		test(64'hdf475b7a25a0aa58, 64'haba316e556927d0c, 64'h00000000b9d61452, 64'h0883040112102c00, 64'h74fda7b50a5285aa);
		test(64'h4e73ad4c42ed9af6, 64'h191a35fbaad63c43, 64'h00000000ada41d36, 64'h010011d982923842, 64'h27ec5b23247b95f6);
		test(64'h4b5a5529ee72e0fb, 64'h2d906c24cafd5bfa, 64'h0000000159bdc43f, 64'h0d806804c0b803ea, 64'hfeb0d8bb86555a1e);
		test(64'h9977f213a8db1fcd, 64'hbff6596f2fd0fab2, 64'h00000165fc0f1c78, 64'h04e4406628d0f0a2, 64'h4f37a27ef84c66dd);
		test(64'h63ea3e237569b7c7, 64'h3c38b203b5c67568, 64'h0000000022bef47c, 64'h3410a200a5466068, 64'h6975c7b7ea63233e);
		test(64'h40482e094a99a382, 64'h6fab817caa9e3045, 64'h0000000080808f90, 64'h2288811880980004, 64'h0848d16058663514);
		test(64'h27b578984885bd65, 64'hf360e0c570694f5f, 64'h000000005ae20b65, 64'h2100400130294545, 64'h191eade4a6bda112);
		test(64'h920d2c369d33aa01, 64'he73b7b2913896d15, 64'h0000000222a92961, 64'ha132312811080001, 64'hc19316e05520e633);
		test(64'h429bf945bb499a8f, 64'h6ca98aa045fc4a7a, 64'h0000000022f05263, 64'h68a102004468403a, 64'h2f6a16ee15f66e18);
		test(64'haf719f4f2bf66c6e, 64'h082a41ab33db5b36, 64'h00000000313df54b, 64'h080841aa30ca0a34, 64'h39b9e89ff6f1fa4d);
		test(64'h73a0e986380ce000, 64'h73f8585358c4f9c0, 64'h000000007e9499e0, 64'h3200180340000000, 64'h73a0e986380ce000);
		test(64'hd65977cb50150033, 64'h42b59a14ee1546f3, 64'h0000000065510e0f, 64'h40800204400000c3, 64'h00cca08aee3db6a9);
		test(64'h23a73d548b3ab0be, 64'hab52c245ee292a5f, 64'h00000000591a5d1e, 64'h81120244a600085e, 64'h2abce5c47d0d5cd1);
		test(64'h6403de97d5620fcb, 64'h13094117519a5914, 64'h00000000000dfc4c, 64'h03000100119a0814, 64'hed794630f0bc5d26);
		test(64'hc3b9596903c1a8a6, 64'h4a8378929056c277, 64'h000000000b6c1116, 64'h0283001210104046, 64'h1565c0839a96c39d);
		test(64'h3440f9dd5cee1233, 64'h62e59bce5a3b22d7, 64'h00000002477dd64b, 64'h4245838e002200c3, 64'h9fbb2c0248cc3a77);
		test(64'h006f30122eb90152, 64'hb9fca6324b2e67d0, 64'h000000000da36c0b, 64'h8174260200022240, 64'h3012006f01522eb9);
		test(64'h1872cb3eb6e5cf1f, 64'h2e24a1e98d9a2341, 64'h000000000254d50d, 64'h2a2401680d802341, 64'h24b1c73d79dacf2f);
		test(64'hfd995bb9b2efe747, 64'hb53cbc0994090949, 64'h0000000003ec6f6d, 64'h951cb80190080049, 64'h66fe76a7df718bdb);
		test(64'hc9d3bd01767c691b, 64'h56ddb9ba08bbb709, 64'h0000000473f01c47, 64'h04d519a008910609, 64'he3c6027ebcb92796);
		test(64'hba91641060e82227, 64'h0a85b21649239ba3, 64'h0000000007524827, 64'h0005900008010223, 64'h6071444ed5986280);
		test(64'h56364982f68b5454, 64'ha8c26d0e94c1d7fc, 64'h0000000006a7d715, 64'ha882480490814150, 64'h4545b86f28946365);
		test(64'h157a7e2dd5c42b53, 64'h2c324f02558517c5, 64'h0000000001fe7e35, 64'h2430040011050505, 64'ha25bdbe1ae8c713a);
		test(64'h266a849f0bc74caa, 64'h584ccc017cf0a8b3, 64'h0000000001a62c3a, 64'h484c040150c08822, 64'h23550d3e129f4665);
		test(64'h34ffd4325d710522, 64'h16a3e6fe9a7eefa8, 64'h0000006fd196e02a, 64'h060246ae02024420, 64'h715d2205ff3432d4);
		test(64'hf11c87d3d5eaf877, 64'h000d9f77f77fd047, 64'h0000000d3d7b757f, 64'h00019a575370d007, 64'h8f38e1cbab571fee);
		test(64'hfc32dd808123de27, 64'h36b2ae1a53a4f05b, 64'h00000000e7b015a3, 64'h2002080a51a4100b, 64'h10bbc4f34eb74c18);
		test(64'h6cfb27cf8ec2cf7b, 64'haf6522bc10c9f425, 64'h000000001cde6ccd, 64'h0e60009800c97405, 64'hd41cfc7bc97fb1fc);
		test(64'h80ec0dc7f90bce8d, 64'hb750c0b4f97bda50, 64'h00000001044fe3ec, 64'hb700800478390a10, 64'h0dc780ecce8df90b);
		test(64'h0851b94fc6fdb9e4, 64'h5d201356260cbb97, 64'h00000000045b7fb4, 64'h0c201352220c1b04, 64'h9df2108a9d2763bf);
		test(64'hdb857e01d05ca720, 64'he9a96ee1fcedd66e, 64'h000000dcfc745a68, 64'h0009480170a1c200, 64'h350708da52e740bd);
		test(64'hb240c68612285642, 64'he2501969320dd66e, 64'h00000000170071f1, 64'h8200084010098404, 64'h28848195018e9293);
		test(64'h6a1276f5f5559642, 64'h871aa3ea22ceedee, 64'h0000000156e4a891, 64'h831a214820c26104, 64'h555f819684a95f9d);
		test(64'h823819670fe7cbb5, 64'h22c3539253b84962, 64'h00000000020a4f3a, 64'h22c3039202b04842, 64'h0fbd3ee528c2469d);
		test(64'hbf8d5b94d2c12170, 64'h6848e04a9166ff32, 64'h000000000d43410e, 64'h4040c00010202e00, 64'h84d078345e61ef27);
		test(64'h16ac3539fe85be4c, 64'ha8d22b41d7bea630, 64'h000000000897e8bc, 64'ha8d0200153b20600, 64'hbe4cfe85353916ac);
		test(64'h274bbb69c186577c, 64'hcc39bca1b0db04d2, 64'h0000000004fce456, 64'h00180c0120d304c0, 64'hee968d1e5dd33429);
		test(64'h59059a6c2957c65b, 64'hf56c370762119f17, 64'h00000000a8aa2e6b, 64'h1108250740018513, 64'h59369aa063da94ea);
		test(64'hf68c7452e88299e9, 64'h32d65881b3fcc69a, 64'h00000000f2c6208a, 64'h324040002264c482, 64'h58d123f9b66628b2);
		test(64'h3c724cd06457d997, 64'h54b7c46dcd93f3e4, 64'h00000006d3829f59, 64'h00148024cd126164, 64'h46759d79c327c40d);
		test(64'hbf2a1035568ead03, 64'h3bf477c06b1a9099, 64'h00000000f90824e1, 64'h12d016804a100009, 64'h3a20157f035e4da9);
		test(64'h70ca9ca1388ba3f8, 64'h2e965e1db9134abf, 64'h000000044b85ccf8, 64'h04160404b1004ab8, 64'h1fc5d11c8539530e);
		test(64'h61441d25e83023ea, 64'h21e2364859cff92d, 64'h00000000d18a009c, 64'h21a000480008f824, 64'h034d5d318829a1e2);
		test(64'hb1f3e0445e998d9f, 64'hf6e01ea8337c3944, 64'h0000000059c0318d, 64'hb6400c2801581944, 64'h1b3f0e44e599d8f9);
		test(64'h1133048e1b501036, 64'h759620a32a487d96, 64'h0000000005553887, 64'h6512000002000514, 64'h10b244cc049ce405);
		test(64'h3222a203606b48ed, 64'h718a215a1f1c053c, 64'h000000000318408b, 64'h00882052040c0434, 64'hde84b606302a2223);
		test(64'h7533f97508e8f236, 64'hcfb8efde1a276e52, 64'h000000156f2d28cb, 64'hc50087421a020c50, 64'hf6d5d5ccf8c902b2);
		test(64'h86602ec62a1ef40e, 64'hb61a64beebba0a66, 64'h0000000261c671c3, 64'h8208401e6a800064, 64'ha8b41fb09209b893);
		test(64'hbe0cd1fc764727f2, 64'h576eceb2d1e6153d, 64'h000000071b1ccb78, 64'h506a841281261524, 64'h1fb1b89bcf2ec0d7);
		test(64'h44ebfb6963c93657, 64'h8e8d11adc67fd1fb, 64'h00000005bb56492b, 64'h0885002d0426c0ab, 64'haec6396c69fd7d22);
		test(64'h9c80284099083098, 64'hce95935d51d706f9, 64'h00000005a020c026, 64'h0414100800c00460, 64'h643004668014406c);
		test(64'hf62d39c1130236b4, 64'h329b1f6828cd1fd9, 64'h00000001cb9802d4, 64'h2011100800491590, 64'hc2361ef978390123);
		test(64'hbd5e2605cf6c53a6, 64'h3cc289f2d090a281, 64'h0000000001ec0306, 64'h2c4200a0d0100280, 64'h7ead190acf9ca359);
		test(64'h39a920d502410384, 64'hd2b0d777d973e083, 64'h00000001602d0444, 64'h9000110100320080, 64'hc95940ba04280c12);
		test(64'he9ccbc53992d4782, 64'hfb6bf995a6a4bd8d, 64'h00000075a5cb0c38, 64'ha34321148404b004, 64'hcc6d3ac7e16614b8);
		test(64'h7ae69935dc1b37b6, 64'hed740dc38f2a2c59, 64'h000000007368f1d4, 64'hcd0005420d2a0c18, 64'h3a66d9b5793b27ec);
		test(64'ha5a8eab61bb64e41, 64'h12a9722676e0929d, 64'h00000000076f2d21, 64'h1229302422c01001, 64'h975d45a528d89772);
		test(64'hf3934777398a54f8, 64'h2c46a4e003517e51, 64'h000000000212d156, 64'h0c00842001103e00, 64'h8bbbf363a8f43645);
		test(64'hdaad6047e91868ed, 64'hdaf48dc5ab35c37c, 64'h0000000fd41fa89b, 64'h5ad0084403104334, 64'hde86819e7406daad);
		test(64'h0a7e0a2bba88f7fa, 64'hddada9fee0155895, 64'h000000008e22b46c, 64'h59a4808ea0155884, 64'h507150dbbf5f5744);
		test(64'hca6c36345d59f764, 64'h9dfb520066661d8a, 64'h0000000028d1d458, 64'h1caa120064641880, 64'h933ac1c9565791fd);
		test(64'ha6b65148dafef331, 64'h854021a0efbfe297, 64'h00000000626afde9, 64'h81400120eeb98281, 64'h8a12656dcf8c5b7f);
		test(64'h2829afba0ceed892, 64'hba12635d5b1561a3, 64'h000000002876114a, 64'h0a0062594a010102, 64'h0377b19441495fd5);
		test(64'h80ca2a310f8f43a0, 64'he3a9dfbe0c7ab527, 64'h000000214298c618, 64'hc0805e1e0402a400, 64'hf0f1c2050153548c);
		test(64'h9df4d2daeb71e98d, 64'ha6f7af722dd0c91e, 64'h0000000af915ebf6, 64'h84e58e122910801a, 64'ha7871f76726b4deb);
		test(64'he18490287a82ef0c, 64'h4beb321d8489a9d2, 64'h00000000260484f0, 64'h4aa0020d048900c0, 64'h6082b421bf03da28);
		test(64'h8ae08228b4d28e01, 64'h24a7de2a96628b5d, 64'h00000000310eebc1, 64'h20a2540880620001, 64'h41140d5420d41e87);
		test(64'h4d225cf17891390b, 64'h10b8391aea7d39b9, 64'h00000000234713e3, 64'h00b8010208382029, 64'h073662b4f2ac118e);
		test(64'hb28f9d3cfcc48d8a, 64'he4e819ff698d2611, 64'h00000000a9e79d48, 64'he4c0182428880410, 64'h6e3c714f4e45fcc8);
		test(64'h5056fa8c60ef981d, 64'h7ee019eb7011e06d, 64'h0000000050b49987, 64'h606011e860000069, 64'hfd09e2469a0ac45f);
		test(64'he72bf00e6f5e78ed, 64'h4b24bf98d5bb5f5c, 64'h00000017702b3b8b, 64'h0b00af10d43a0e54, 64'he00fb27ede87e5f6);
		test(64'hc9a5c83d1ce87ee2, 64'h2ead8953fe2c569f, 64'h00000004de51dbe2, 64'h2a058052862c4682, 64'hbc13a593477e1738);
		test(64'h6c4e4957cbf249f2, 64'h56bddadaf20b91e1, 64'h000000050ca6e51e, 64'h5689da1090039120, 64'hc7f186f19c8d86ab);
		test(64'h7f1827fd0a33de82, 64'he87c47b6b47e59bf, 64'h000000399fc0cf42, 64'he850028284765102, 64'h417bcc50bfe418fe);
		test(64'h687d9f75582f2acc, 64'hfe14aa00d33e4799, 64'h0000000034ed972a, 64'hb0008a00c1144490, 64'hba6fbe94cc151fa4);
		test(64'h598db2f22f56fd56, 64'h4fe1d2cd4b45c52c, 64'h00000000ccde1f79, 64'h05e090c54b048428, 64'h65f265dfd8952f2b);
		test(64'h63f67b5db34b85a6, 64'h4099a25fdc22bb2d, 64'h0000000071fb461a, 64'h0090a045c002320c, 64'h783795a49f39ea7b);
		test(64'h8eeb85cb1667951b, 64'h7a3d94d312ef7cf1, 64'h00000003addedca3, 64'h2a04905012c520d1, 64'h6a27299b4ac74dd7);
		test(64'hbbf178749c1bbe48, 64'hbd961c2a326d1b34, 64'h000000007b9a22f0, 64'h1c00182a12681100, 64'heb84c9b18747bb1f);
		test(64'h8749c080462d8c02, 64'h498d83505376979a, 64'h000000000ac29541, 64'h0088025012140008, 64'h2030162d08238719);
		test(64'h744dbf2144ecdc35, 64'h4b09893af74ea8cd, 64'h000000008fc24ea3, 64'h0801013295480889, 64'he88b21f7cd88a3ce);
		test(64'h6e23825bc9aba6dc, 64'h4b64ea8ded28c691, 64'h00000000728aebde, 64'h4104a20d45088680, 64'h41a79d1359ecc657);
		test(64'hac9475a482a9135c, 64'h6a10233c6f77167a, 64'h000000006d9091b6, 64'h4000022844230470, 64'h534ca628a1d561a3);
		test(64'hedb510c9650f26d6, 64'h8713c5bccae04d1b, 64'h000000006d09202a, 64'h841100b840c0490a, 64'h3980da7bb6460f6a);
		test(64'hd6e911d25447ab41, 64'h0ee2d537bcc3d457, 64'h00000003e2a8af11, 64'h04424021b4419001, 64'h884b6b97d5822ae2);
		test(64'h01399961d5bba63f, 64'h235390ec7158beb3, 64'h000000002bb2de6f, 64'h224290687040a2b3, 64'h56cfbadd996808c9);
		test(64'h5419527d6e5fc30e, 64'hda39a46d05027f08, 64'h000000000638fd87, 64'hd029a46001020700, 64'h19547d525f6e0ec3);
		test(64'h36e0cc29a39ab9f6, 64'h486fb13023473105, 64'h0000000000c22e5e, 64'h4846903020472104, 64'h930dcc613556679f);
		test(64'hf351cfe8c8a35e27, 64'hd59b3b13b897715b, 64'h0000000ea4e26743, 64'h81820900a817010b, 64'h713fa8fc4ea75c31);
		test(64'hceae16bb86e36979, 64'h2537dc9c87cdd1eb, 64'h0000000562f7655d, 64'h2130549006c441e1, 64'h7c16e9695737dd86);
		test(64'hd6e2ebeb569b5088, 64'hf6fc27dcc4a14429, 64'h00000000df8bd3b2, 64'h52a4234800800400, 64'h67a944a0d1e9d7d7);
		test(64'h128f4bce243e2ce1, 64'h3eaf8695e39148f8, 64'h000000009bcd113c, 64'h0420869043014808, 64'he12c3e24ce4b8f12);
		test(64'h4ec5caa4adc95469, 64'h0d3905364548fc81, 64'h0000000003094f55, 64'h0521002441006801, 64'h8dcac5585ec6a896);
		test(64'hc9cc3adebe1d6d38, 64'hcb8491fd1a5919e2, 64'h00000000775bbbb2, 64'h4b8000e912480980, 64'heb4797c23633ca7b);
		test(64'hd0aeeefc73b59351, 64'h09fc2af3cc320c37, 64'h0000000015ff1309, 64'h099c0a5240300821, 64'hc98acead773f0b75);
		test(64'ha21dda8c6d7185ef, 64'h8666fd63e33ffd24, 64'h000000296c06e30f, 64'h0240d9230302f524, 64'hd61758fe2ad1adc8);
		test(64'h71753d42831e4bde, 64'h7886c619896340c9, 64'h0000000003910a5e, 64'h6006c010816240c8, 64'hbab2813e2d43ed87);
		test(64'h58b269aaa2a89408, 64'h72a4ad17c109c720, 64'h00000000056694a8, 64'h2220810280000400, 64'ha2a8940858b269aa);
		test(64'h55f171a0ad421cae, 64'ha6b310d419247317, 64'h0000000002ee1846, 64'ha220008009202216, 64'h8e05aa8f3875b542);
		test(64'h448e2c074a0a1e31, 64'h3195d373c945a64d, 64'h000000001401b031, 64'h1011005009440601, 64'hd488b0c1505823d2);
		test(64'h30f3cbe1f7f51e41, 64'h9cf63fdfe2ef443d, 64'h0000009e9787faa1, 64'h9c063bdd406c4001, 64'h28d2afbf2d7c3f03);
		test(64'hebb1c4fd659635f5, 64'hbbb64c42b5d2c4de, 64'h000000037e59767a, 64'h2a2604028190c4ca, 64'h7f134eeb5f5c9659);
		test(64'hbf405fea313d96d7, 64'h7228523f6894b83a, 64'h000000000e7a93a5, 64'h402012362090a81a, 64'h7d69c7c4ba5f10ef);
		test(64'hb838288a1bf8dfca, 64'hce16ed21d3eb9cf5, 64'h000000148607f3f0, 64'h4400cd21c0cb9c24, 64'hfe5c724f41544743);
		test(64'h76718099b42dd68c, 64'ha00e1eb36aa3ae21, 64'h00000000080aa2cc, 64'h800804a348a10600, 64'h781ee94cb9b24066);
		test(64'he51e61b25323413d, 64'hde795564468ce8ff, 64'h0000000c8d2a843d, 64'h122141004480083d, 64'hbc82c4ca4d8678a7);
		test(64'h19211646edf82eee, 64'h0b422f855193a533, 64'h000000000a195c6a, 64'h0a422e001092a432, 64'h47777bf186268948);
		test(64'h8f577643160daeb9, 64'h340b6791d1d53ba4, 64'h0000000017e243b6, 64'h04030090c1542b04, 64'h61d0ea9bf8756734);
		test(64'h0668ef89d1eaf8d3, 64'hd79129c5142979e2, 64'h00000000061e6ded, 64'h4191088514203122, 64'h74baf27c0992bf26);
		test(64'h43e1ae909c411391, 64'hc21ac4fc24a355f6, 64'h0000000031644564, 64'h0218040400205442, 64'hc4463641ba06c14b);
		test(64'h0e6177ebc33baedd, 64'h4ffa6888320dcec0, 64'h000000000e6366df, 64'h0338680812098e40, 64'h0e6177ebc33baedd);
		test(64'h72c68990d278655d, 64'h5743b824a4c062d7, 64'h000000000d69239d, 64'h0443800480804255, 64'h91094e63a6ba4b1e);
		test(64'h65cc0172be6fb7d2, 64'hc00dfe1b8e7edc3d, 64'h0000000700afdea8, 64'h00097c0a8e5ad824, 64'h1eb7f9d71b20cca9);
		test(64'h5aa6e86ee0d88ec5, 64'h429e57d947d22e98, 64'h00000000e705473c, 64'h4280158101c22088, 64'h6ee8a65ac58ed8e0);
		test(64'he2cf3dd71d8f2cc5, 64'h6ecb5e15725fa3dc, 64'h00000019fbb91e99, 64'h4e034c0170162214, 64'h7dd3fc2e5cc2f8d1);
		test(64'hc27f95eeec1e6b9b, 64'ha9583aa25837d18c, 64'h0000000011d3d72e, 64'h28001a805027110c, 64'hf72cee59e1ceb9b6);
		test(64'h7ddfbfc3511c5d2f, 64'hbfa5ac5287a6ce55, 64'h00000003dbfa24e3, 64'h3501045002a48455, 64'hf73cebfeeaf12ac2);
		test(64'h4c8586fe7fc2b689, 64'h068ab7174609b1a4, 64'h000000000526ee74, 64'h068a021306010104, 64'hf72c6b98c45868ef);
		test(64'h4e1b36d34b534bc7, 64'h929c7dd9a94ffc90, 64'h0000000166ba734a, 64'h12105941880bc490, 64'h36d34e1b4bc74b53);
		test(64'h11de6a8138a24769, 64'h7f2be451a9e1f9a7, 64'h00000004598b5229, 64'h042a20402080e921, 64'h1c45e296887b5681);
		test(64'h2638093e2ad0b394, 64'hc0a81a4a1b3d77f3, 64'h000000001a6c86e4, 64'h0088084810151650, 64'hdc9245b009c746c1);
		test(64'hf55946cecd1091dc, 64'he09f9378896b47ff, 64'h0000001d929e01dc, 64'h608c9108002101dc, 64'h3b8908b373629aaf);
		test(64'hd477f7fe57378eb0, 64'h7018023a0cf64dad, 64'h0000000005be9ed8, 64'h7000022a0c160980, 64'hb3ba07d4bb8edfbf);
		test(64'h8af8e4b158256a76, 64'hb3172f2864c57d22, 64'h000000004a2943d3, 64'h9200222060843920, 64'h52859ad92af2b1e4);
		test(64'hd9b092185447ff58, 64'h35276a56c7b7a6a6, 64'h00000002c0a307f0, 64'h00224040c7b72280, 64'h15d1ff25670e8624);
		test(64'h0a578fce33d3a06b, 64'hd0174b85d4877deb, 64'h000000007be2b41f, 64'h80060b81148201a3, 64'hbccc6d50ae05371f);
		test(64'h44fb1c6fc2ec69d0, 64'h34cc5f69a14fc503, 64'h000000001e73e714, 64'h20085b0181074000, 64'h22fd836f347369b0);
		test(64'hed729b2e2dce7a49, 64'h5f3eeaae64b854fd, 64'h0000002dccdee725, 64'h4e0aaa0e04b04091, 64'h685bdce1d1761bed);
		test(64'h6385c9826ad3bb14, 64'h04a3b4c51f4e5962, 64'h00000000098854b8, 64'h0082a405170c0840, 64'h9a7cee419c253628);
		test(64'hb0da7a97376add50, 64'he4f2bd7021cd5cea, 64'h00000002b6e1d9e8, 64'hc0d29920214c4880, 64'h9acd50777ae06dda);
		test(64'hb24c32b260e2bcd3, 64'ha0d49c7f31c22d6a, 64'h000000006a8ca7e9, 64'ha0001c0a3180290a, 64'hb8907ce313e8e8c8);
		test(64'haa5a39bc9de7b3b0, 64'h0e1fa7d94ae890d7, 64'h00000001749b2ee8, 64'h040ea6590a2880c0, 64'h9c3d555acd0db9e7);
		test(64'h7423e71e782f9436, 64'h5846d333b080069e, 64'h00000000031db34b, 64'h0004d3028000028c, 64'hb4dbc81d9c16f82d);
		test(64'h4bf70a0f35156113, 64'ha90a057e1c276f11, 64'h000000000683d5c7, 64'h8808005418010411, 64'h050f87fb92233a2a);
		test(64'hf298853a8f38c58f, 64'hb513f238432e37c4, 64'h000000007243bc2d, 64'h05127008400a21c4, 64'h2f8958a3f8835cf8);
		test(64'h6d902e130b8b1aab, 64'hbf7bb3e320b3c65e, 64'h0000001690a1a625, 64'h2609a0a200314216, 64'hc4b80679eaa4e2e0);
		test(64'h7820bdcb5e6cf652, 64'ha4137fe53b5bfb3e, 64'h00000041ee5d4f49, 64'ha0026bc12a1b6224, 64'h859f39b5e37e082d);
		test(64'hc406b657de244348, 64'hb8f934cbc37dd9ce, 64'h000000200ebe492c, 64'h28f134024020c840, 64'h9013d59e18b721c1);
		test(64'h8726ed54134e91fd, 64'hb5fe02041dcfd39e, 64'h0000000264d97abe, 64'h009a00001c84539a, 64'h157b98d27f46b1c4);
		test(64'h8c28c4584b016bb9, 64'h80cea7d758e6a72e, 64'h000000024a3140bc, 64'h0008860048a2a322, 64'h40e16ee928322513);
		test(64'h1c381264d8db61e0, 64'hde92f77015c8af23, 64'h00000000e42b4e8c, 64'h1a8066601400ac00, 64'hb1bd687083c18462);
		test(64'h9939287bbf5696bd, 64'hdb12ad9a26fa34d0, 64'h00000000b663f55d, 64'h9b12249202683490, 64'h287b993996bdbf56);
		test(64'hda937fd603d2f4b9, 64'h6da5672dbbdf5f10, 64'h000000293f20f969, 64'h2500032913c91c10, 64'h7fd6da93f4b903d2);
		test(64'h632fa8ccb7c125ae, 64'h338ba6ece2980c65, 64'h000000002df37716, 64'h318b004420900864, 64'hb72ca1d539f145cc);
		test(64'h6a4daf6f96a8853d, 64'he41cfb0785ed3b77, 64'h0000000cebfd605d, 64'h6418590280402875, 64'ha1bc6915f5f656b2);
		test(64'h9cd05e20ef44dcc1, 64'h40a5a3256e454538, 64'h0000000001053fb0, 64'h408402052c050008, 64'hc1dc44ef205ed09c);
		test(64'hecc8b62f1e0b81b2, 64'h65722a86c683ba31, 64'h000000001d159b86, 64'h6500088600019810, 64'h42712d07791fdcc4);
		test(64'h4f068efe3eac1105, 64'h68972c52bb3ba867, 64'h000000014cfbd405, 64'h0097084280210005, 64'h7c3588a0f260717f);
		test(64'h0f800a95e84526f7, 64'h2b2bfef794f6f17a, 64'h000000e0166c489d, 64'h0822f4108422b15a, 64'hfd8915b2650a200f);
		test(64'h98bfd6e99c7c0218, 64'h23ff80a2283f7c1c, 64'h000000000bfe7c06, 64'h01c7808000020c00, 64'h9e6dfb898120c7c9);
		test(64'hf6110a4987fb85e4, 64'hc371bf908d778bef, 64'h00000038c517dcf4, 64'h02300f90896083c4, 64'hdfe127a1886f9250);
		test(64'ha7aea886fe827f38, 64'h652b33b7778bb5c6, 64'h0000000fd137d4f0, 64'h050b3320238b8580, 64'hdaba2a92bf82fd2c);
		test(64'hcea27c9eab6b132d, 64'h15739799720aae4b, 64'h000000004a672e15, 64'h1123151810028449, 64'h543797e36d5d4b8c);
		test(64'h161897b3042249d7, 64'h51556ddc128a9884, 64'h000000000241d027, 64'h4004088802888884, 64'h6181793b4022947d);
		test(64'h99b3846002732cb5, 64'h1ea18d72b47247ac, 64'h0000000067ac0f4d, 64'h00200d1210604324, 64'h37205bc23b990648);
		test(64'ha7c7ceb69538c823, 64'h22fe60600dc2d173, 64'h000000000f1cb18b, 64'h024e002008800103, 64'h314c9ac137d65e3e);
		test(64'he5184b9d37616811, 64'h98e4ca04e5558e81, 64'h0000000004079e51, 64'h98600200c4000801, 64'hda24876e3b929422);
		test(64'h3da10e5a4394a5dc, 64'h391b9fa671af7b97, 64'h000000789c33223c, 64'h290881a050245a94, 64'h705abc85a53bc229);
		test(64'h541bfcf0f8a020a0, 64'hfb9482b9a48f48e1, 64'h000000002857340a, 64'hf084000080024000, 64'hf4501050a827fcf0);
		test(64'h099c0b5481684e30, 64'h657981315ee712ac, 64'h0000000009940614, 64'h0011802008e01200, 64'h861803e4c99045b0);
		test(64'h7e85da2f88d9f789, 64'h928e15ebd3088626, 64'h000000000750f878, 64'h800c146b53000202, 64'h2267df62bd52a7f8);
		test(64'h4238a5c26b1fdeaa, 64'h84cc4ea6c4c50b97, 64'h000000000114a3d2, 64'h044806a684c40912, 64'ha543421c7b55d6f8);
		test(64'h432695eb11fc8440, 64'h10ce90d7f2e66d48, 64'h0000000007e62f0a, 64'h004090d640404000, 64'h2643eb95fc114084);
		test(64'h4ffd9435ce15f392, 64'h4bd8e6a2676d7cf5, 64'h0000001ff2561f24, 64'h42d06400456c3844, 64'h3f16dca286a3f8ef);
		test(64'h31941ddf21fa3b4c, 64'hff6ceaae9e2a9c3a, 64'h0000000c44570762, 64'h7c406aa40e0a1030, 64'h13cefa847f4761c4);
		test(64'hf4cf7f7415328782, 64'h67447cbb6553420d, 64'h0000000073fb06c8, 64'h0504182805500004, 64'hfc8f8bfb13a214b4);
		test(64'h8560e820a09ac7c9, 64'hf2c30aeddf9f2006, 64'h00000001048881d0, 64'h50000864c3990002, 64'h52092b080aa6d363);
		test(64'h8a4183adb864dfc6, 64'h02d09f7e2e2927f9, 64'h0000000151ad91f0, 64'h029090640c292718, 64'hc9ef98745e438245);
		test(64'h5901dd892b2fabf6, 64'h504f96c695afc921, 64'h0000000061e817ee, 64'h100b04c6848fc120, 64'h171f57f9a602ee46);
		test(64'h76257e5e77b4fef3, 64'h03ce1ebd2e264bce, 64'h000000010bcebdd9, 64'h00ca1ca82e260b86, 64'h589db5bd1eddcfbf);
		test(64'hd187a12d7d2334d9, 64'hb0c1598ac06f64f0, 64'h000000000b4529bd, 64'ha080408840494490, 64'h34d97d23a12dd187);
		test(64'h59cfa4d52eda8639, 64'hfa176ecf580b9d75, 64'h0000000b3ab53a4d, 64'ha805664a40018161, 64'h9463d15e85ae6afc);
		test(64'h266a772159ec770f, 64'he9169de3f6e18c21, 64'h0000000042b2a9c5, 64'ha1109cc0e6800c21, 64'ha6dcbb0f1995bb12);
		test(64'h572cc72f76196779, 64'hb929bf38d5adabf7, 64'h0000002e8f5c55b9, 64'h11293b00508c2af1, 64'he69e6e98e3f4ea34);
		test(64'hfe5fcce3a0d2ed60, 64'h78dc22802ff010ba, 64'h0000000007bcc348, 64'h089020802b501000, 64'h90b778a0bc335ffb);
		test(64'h83149c49ed8a9e1b, 64'h25ca04d194fb6de7, 64'h0000000042b63183, 64'h258a00c010a36063, 64'hb75179d8c1283992);
		test(64'h49de5f48614d02fc, 64'hf8bd38e64d62a7f9, 64'h00000009b9a260be, 64'h40301086080023f0, 64'hfc018e9284afed86);
		test(64'h3a4fa9f5f442bcf6, 64'h24494464d085c40f, 64'h00000000005cfc56, 64'h20004044d001c406, 64'hf25caf95422f6f3d);
		test(64'ha74d5460d85a2c47, 64'h96305827995769df, 64'h00000001668ed327, 64'h1430000588054087, 64'h062ab2e5e2345a1b);
		test(64'h18b81f53cf1c50cc, 64'h9f9e89629355db6d, 64'h0000000638edb316, 64'h0f0e802280440a28, 64'hc2fccc0a47423af2);
		test(64'h3353ce6e2f5e0b9b, 64'h252efc708769314c, 64'h0000000028e79e8a, 64'h212cbc000268110c, 64'h3533e6ece5f2b9b0);
		test(64'ha1dc9940fa5e302e, 64'hec9f3b41a5bf47ce, 64'h00000029e36c3c07, 64'h001f1101a418014c, 64'h374a0166b5afb80c);
		test(64'hc833a251b45e0ac1, 64'h72e6e42b8cc42694, 64'h00000000105a1acc, 64'h5022e00084440004, 64'h2a158c33a01c4be5);
		test(64'h0a0f8e9579b48bd9, 64'hcdebc5dcc602348e, 64'h0000000020f5540c, 64'h4d29844086022482, 64'hf0a056b21e6d67e2);
		test(64'h4f778e831f5cd367, 64'hfabe0ac6f2385301, 64'h0000000026df237f, 64'h3a96084492180301, 64'h8fbb4d432face39b);
		test(64'h09c0ee797c66c3e7, 64'ha8cb40d2601217a0, 64'h00000000001c5b4f, 64'ha0494000601211a0, 64'h7c66c3e709c0ee79);
		test(64'h9cc3ab8e35bddb8f, 64'hfba6f240ba21a3f8, 64'h00000001326a6771, 64'h1924f040aa01a078, 64'h8fdbbd358eabc39c);
		test(64'h5438364aba3c1ebf, 64'h55cac4ff711c2942, 64'h000000007114a6e9, 64'h154044c170142942, 64'h51c2c91aeac34bef);
		test(64'h0c5d1b314efc0190, 64'h2773622c28759d93, 64'h00000000254c7c1c, 64'h2163622000009100, 64'h8dc803ab089027f3);
		test(64'h5e79370c3a207268, 64'h7a38c923f51da88c, 64'h000000005f883012, 64'h3820400070118800, 64'h97e5c07302a38627);
		test(64'h7e040ff7213630dd, 64'hc20997c1d31bcbfc, 64'h00000000c3f0d037, 64'h80080241500a0374, 64'hdd0363127ff040e7);
		test(64'h6ce39098e9e6836b, 64'hc7b38f4e98a2f4ad, 64'h000000033704be0d, 64'h03908e0c8000d425, 64'h9d6d79343dc94606);
		test(64'h66f20f9407b33a04, 64'h3bb7c6181ed25d70, 64'h000000012e8e3b60, 64'h0036c01806900040, 64'h3a0407b30f9466f2);
		test(64'h9a618fe49a42a5ca, 64'he7e10859b3641201, 64'h000000000227c5a0, 64'h8420081093040200, 64'h65924fd865815ac5);
		test(64'h13f55cc5af8c7a65, 64'hdcd1a3e4ff235bd1, 64'h00000004f0daf1e5, 64'h1490a380c7210a41, 64'hacca23fab59a5f4c);
		test(64'h258d4c9b073dc926, 64'had4e9eee310d3b34, 64'h000000016c694f2d, 64'ha00686ce01010830, 64'h9c6270d3c4b952d8);
		test(64'h82926cf0d1c36c42, 64'h12d834425907ba1a, 64'h0000000001ab6b51, 64'h02c0044051042008, 64'hf093682818933c74);
		test(64'hab4009ac8cc473ee, 64'h4d29a67debaec089, 64'h00000000a016924e, 64'h0809060868ae4088, 64'h80575c06c84cddb3);
		test(64'hd769908f1d489f48, 64'he33206b9fa50dc76, 64'h00000001b84c6af0, 64'h813004882250c820, 64'hf621742106f2d769);
		test(64'h45a2ffbb4681a04e, 64'h62ea749f4571708e, 64'h0000000095fef0a7, 64'h202840064000408c, 64'h8a51eeff4291b10a);
		test(64'hf2337c65ea6871ef, 64'he1d1d590c0053acc, 64'h00000000071b8ccf, 64'h40c10190000138cc, 64'h332f56c786aefe17);
		test(64'hcec3852f40e003b9, 64'hfcc8edc53dea0dfe, 64'h00000067a33070dc, 64'h5c8800c400000d72, 64'h6ec00b01f852c3b3);
		test(64'hb56bb3b640676665, 64'h4000f2a8fa2091e9, 64'h00000000005f210d, 64'h0000c2a0ca001121, 64'h9b809a99977a7973);
		test(64'hd28725ac24d98a8a, 64'hbeb43332cd9ddb1f, 64'h000000299982ecca, 64'h98101030c181480a, 64'h35a4e14b51519b24);
		test(64'ha40b2673fac1c769, 64'h6677f8c8e8e6bea7, 64'h00000018322fc469, 64'h6077a88008c0b621, 64'h5f83e39625d064ce);
		test(64'he8631687e3783a1a, 64'h91dce6db2c2f0cee, 64'h0000000440e39885, 64'h91d062d0042a0064, 64'h2dcba4acc92bd294);
		test(64'h15ad6c0b22c7a977, 64'h19dab0ce478c9be5, 64'h00000001648a56af, 64'h10823006450813a5, 64'h11bc65bba2e5c970);
		test(64'hb2c3a87c1c7ddb92, 64'ha10b3327490b84a5, 64'h000000000338c568, 64'h000b3125410a0404, 64'hc2eb7e16173c45cb);
		test(64'hcd856e6a00341aec, 64'h1ce80aeec9dd49d9, 64'h00000000e3740a5a, 64'h0000002a00544950, 64'h959d4acedc253800);
		test(64'h6d6b2c3d8033a50a, 64'h82fa43f402fbc0c0, 64'h0000000001b071b8, 64'h000a01d000a08080, 64'h6d6b2c3d8033a50a);
		test(64'h5f49920022940741, 64'h672f8b0fb926df0f, 64'h000000174d021071, 64'h000409028000d401, 64'h92fa0049294482e0);
		test(64'h56c488d656e0b171, 64'h3b4d56104ce90c53, 64'h0000000005506f0d, 64'h1948020048210c01, 64'h11b6a632d8e8a670);
		test(64'h12c8ae4122afaa8b, 64'h110f77a2906d371e, 64'h0000000050b01f25, 64'h010125a280491016, 64'h41ba2384e2aafa88);
		test(64'h59cc0223bd03eaf0, 64'h12eaead265975125, 64'h000000005a08b8e4, 64'h02e2005261135000, 64'he7305d0f6acc1031);
		test(64'hc1775a75632296c7, 64'h2197a2ce17cd822a, 64'h000000000bca8c19, 64'h00148044058c002a, 64'h889c3d69dd34d55a);
		test(64'h2d8a6d786f9bd3ae, 64'h34712dc19cd7cf89, 64'h0000000143d1d79e, 64'h04512c411c91c588, 64'h451eb49e679f5de3);
		test(64'h09252bbe9740a256, 64'h144200bcc3287692, 64'h000000000007ec4b, 64'h1000000880202490, 64'h8eeb0685a8596d10);
		test(64'h332dcf2bfb9fc2ff, 64'hc9ac46b7f6b3a2ba, 64'h000000017e9fb7bf, 64'h89ac42a3f402a2ba, 64'hff386ffe8e3f87cc);
		test(64'hdbdaced3171f2b7f, 64'hd9d58a40c6462ae9, 64'h000000001fe79bef, 64'h99058a0042060ae9, 64'h2f2bbf17e5e7e3cd);
		test(64'h3b168f976ae53cfc, 64'hbf2d1fcec9ea4985, 64'h0000000764f9b716, 64'h3b090e44498a4980, 64'h7392f4b659adc3cf);
		test(64'hc211a0c8df775c56, 64'ha3445b78b648676e, 64'h00000000a0137a93, 64'ha14453589248024c, 64'hddf795354483230a);
		test(64'h1e2ea88b0190ec20, 64'ha4f96b71e5dcc5f8, 64'h00000004a60869c4, 64'h20c0031005980100, 64'h20ec90018ba82e1e);
		test(64'h7a4faa57ed7f0273, 64'h34b4a701fc4500b7, 64'h000000000c3af7db, 64'h3094a700040100a3, 64'h40ceb7fe55ea5ef2);
		test(64'hc264ac6ec0074776, 64'h1a4b4ff65c485478, 64'h000000001863705e, 64'h100000e40c405430, 64'h764707c06eac64c2);
		test(64'hadbdbfa21dcadad0, 64'hc5bb8fd886d7fb65, 64'h0000005fbf8596e8, 64'h40208dc082535900, 64'he25c5e0ee5e7f715);
		test(64'h8950e4ac26ee2dd3, 64'h418ceb94ca02e548, 64'h00000000011c519e, 64'h408c6810c202a048, 64'h5089ace4ee26d32d);
		test(64'hc125f13c5a82b282, 64'h82cdd70e7a055767, 64'h000000010f9d7142, 64'h008c90022a004402, 64'h5a414d4183a48f3c);
		test(64'hb8a0daee855a6409, 64'h421874c0a74af281, 64'h000000000015d7b1, 64'h40106400a1001001, 64'h7450e5dd4aa59806);
		test(64'h8dca353864a0e724, 64'h0d45a2b6ff60efea, 64'h0000000f13191ee4, 64'h0801808483406920, 64'ha09181bd3a27c2c5);
		test(64'h0f21f5117e3294b5, 64'h8b25d8987b457cdc, 64'h00000000f797c0b5, 64'h8325809028411494, 64'h115f12f05b4923e7);
		test(64'h44e8d0b1b73d4125, 64'h69767dd516e9d2e7, 64'h0000002314579d0d, 64'h60325c5504804085, 64'hedbc82a422170b8d);
		test(64'h2aed3f6e8de85882, 64'h5206ace5f093e8b3, 64'h0000000019dd10b2, 64'h00062ca020904002, 64'ha1141b71cf67457b);
		test(64'hcb31e3ef65da83a2, 64'hd837acc1a18f9e25, 64'h00000000dce77a8c, 64'h50138c4080038804, 64'ha95e34157c233dfd);
		test(64'ha277a21ee25da859, 64'h7bcbed59b76a2549, 64'h000000092e86caa7, 64'h79c0895192020501, 64'hbb512d51aed1a654);
		test(64'h326b2e4a9ca28343, 64'h2547db839c597685, 64'h000000009632f009, 64'h2046480280092005, 64'h1379d158c6153438);
		test(64'h513a808129bcc528, 64'he0d3480a313ff6a2, 64'h000000001182f992, 64'ha012480a01229200, 64'h86e3358254ca2024);
		test(64'hdca282d957ea61cf, 64'h3b08fcbc1e7c26cc, 64'h00000000c416bd4f, 64'h2900fc280c0c20cc, 64'h2acd9d28ae75fc16);
		test(64'ha7ccbaaca692ed81, 64'h08bc118b16e0881a, 64'h0000000000276398, 64'h0024018912800002, 64'ha3ea33ad24b768a9);
		test(64'h58fb3a69b6f80f8a, 64'hfe96d461604d5d15, 64'h0000000059a5dc38, 64'hb616c000004d4104, 64'h53694a7ff054974f);
		test(64'hbf62f9685fa622ef, 64'h3b7c28e1c818356a, 64'h000000001fc6cc8f, 64'h3b5028010010346a, 64'ha95fbf8898ef92f6);
		test(64'h1c9ec79134281f80, 64'hb44807b940c9afbf, 64'h0000000037d447c0, 64'h140800280000af00, 64'h01f8142c89e37938);
		test(64'h16283a5753943320, 64'h3a4b293238d7d346, 64'h000000002a66ac38, 64'h280b011000c31000, 64'h9428acd5c516cc08);
		test(64'h363a928049fa6d60, 64'hf9b2ba35f92ac1ba, 64'h000000031ea09f68, 64'h01103a3131224100, 64'h9097fa162068cac9);
		test(64'h759ceda5f52dbab9, 64'heeb4865a9de66f8c, 64'h00000006af06ccd6, 64'h4ea404128ce22704, 64'hc9575aded25f9bab);
		test(64'h2a1813221c11c053, 64'h782e60a64a759713, 64'h0000000015054587, 64'h3800200248001203, 64'h8c44458130ac8388);
		test(64'h0c248e76989cd8fd, 64'h8f6e1ad7359c7e0c, 64'h0000000314de4fb3, 64'h8a28085431807e04, 64'h42c067e8c989df8d);
		test(64'h679473cef8c945f0, 64'h072288212921ab7b, 64'h0000000001c0c878, 64'h0300800108008b60, 64'hf02a39f137ec926e);
		test(64'h9634ccb3bbac56ed, 64'hf2de849797131500, 64'h00000000132bdec6, 64'hd296001293111100, 64'h9634ccb3bbac56ed);
		test(64'hff3ad229f80c732a, 64'h81d15ff9e41de14c, 64'h000000019645f33a, 64'h81d10060e00c4108, 64'ha3ff922dc08fa237);
		test(64'hd40366b4bf98098e, 64'h0cee390c05ee9a1d, 64'h000000001061e426, 64'h0cec18000022801c, 64'h8799308ed46046f7);
		test(64'h87dd4cc275d26069, 64'h3ee01b25347efee9, 64'h00000001e41e960f, 64'h08e00924204c0641, 64'he1ba9690ee4bc18c);
		test(64'h545cc8388cdc9954, 64'h10e1dd83b305f566, 64'h0000000053410a5a, 64'h0021198221045120, 64'h323766151535232c);
		test(64'h3a6e9fd005aa670c, 64'h84f0b1e9625d70c2, 64'h00000000035e0130, 64'h00b0214140581080, 64'hca9b6f7005aa9d03);
		test(64'h9edb1522fc9bbaa3, 64'h95ce659462f44516, 64'h000000003ba63481, 64'h9508619062504006, 64'h5488b6e7aeca3fe6);
		test(64'h79fcef1d2fba281c, 64'h0d2808a608f4db4c, 64'h0000000001796c23, 64'h0c28082000a00340, 64'hcf97d1feabf2c182);
		test(64'h6c73755f214e61fa, 64'h4275210387d9c3b9, 64'h00000000177c54be, 64'h001100038180c3a8, 64'hf5928d12afbab39c);
		test(64'h112f66f8322dbe7e, 64'hfcf27daf8bedba82, 64'h00000010b97047fd, 64'hf802482689e8ba80, 64'h448f99f2c887ebdb);
		test(64'hb5b632429a2a8177, 64'h489216e516fa69b5, 64'h000000001ea2962f, 64'h0090104412004995, 64'h24bb56511318a797);
		test(64'h58fe77a48f375026, 64'h703b307d0ff5f706, 64'h00000005f6979ea3, 64'h4021304c0ea01104, 64'h25bfdd1af2dc0598);
		test(64'he759944e8ca71d68, 64'h1ed852f9c9700952, 64'h0000000006e92a5c, 64'h0c4802c1c1300100, 64'h611bbd56479223ad);
		test(64'hdeaeaa959c4afdc0, 64'hc9b615c4ca03183b, 64'h000000000ed8b560, 64'hc02204c4c8031000, 64'h30fb25939a5557b7);
		test(64'h2823d13141c070cb, 64'hb75748761892a2ea, 64'h000000002039845b, 64'h805400061000a04a, 64'h30143ed08c82c474);
		test(64'h2e0030de7e087d2f, 64'hb989567cc364c615, 64'h000000002825d833, 64'hb9800204c3204215, 64'h03ded100ebf1db40);
		test(64'h1578b5ae2ea32ad9, 64'hd6ff94454af7facc, 64'h00000019e3a74cbe, 64'h468b84040292b284, 64'h8751ea5b3ae29da2);
		test(64'h82fcd6ebceb72639, 64'hc0d74c2a9c4ee635, 64'h000000005e5f667d, 64'h80550c0a84060621, 64'h9163dcb79e7d14cf);
		test(64'h5e38b78eab7b56b9, 64'ha810f47a5e872e54, 64'h000000000ee3299a, 64'h8800d46a14850e04, 64'h7be8e583659bbab7);
		test(64'hb6595ca3842b3508, 64'hf00be8e0ed8b2162, 64'h000000001756c4f8, 64'h2000a0c064800100, 64'h218ec502e95653ac);
		test(64'h397b8fd375f42fa0, 64'h8d4eb56f741e2fff, 64'h0000005d9c7f5fa0, 64'h8906344f50020fa0, 64'h05f42faecbf1de9c);
		test(64'h61e24c5f70420c60, 64'hca1e4e48bf5d9078, 64'h0000000041ed840c, 64'h4a00080081418000, 64'h600c42705f4ce261);
		test(64'hedf0618021f83558, 64'h2aeb574f7f799332, 64'h0000003711021f2a, 64'h0001014f03288300, 64'hc55284f29420b7f0);
		test(64'h3b20a6dad4adec94, 64'h38cbe46dd377124d, 64'h0000000382e9c542, 64'h2889204cd2620208, 64'h01735e95e58e86cd);
		test(64'he1b0bc06a90ecf29, 64'he43675e14fe438f7, 64'h0000000ec7024491, 64'h602444014b243051, 64'hf39495703d60870d);
		test(64'hbb94ae73a9e72d46, 64'hf3f5cb5737ef729c, 64'h000002f9adb8f741, 64'h93348856164d2018, 64'h37ea49bb64d27e9a);
		test(64'h6de90bee9afd8b79, 64'hae0d628b559b8e2f, 64'h00000000ea793bb9, 64'h2209228b14098629, 64'hbf599ed197b677d0);
		test(64'h62081805f1f0d2f3, 64'h0f258f844355ef96, 64'h000000002086e62d, 64'h0f008f0001444f06, 64'h2450892087cf4f0f);
		test(64'he46aeb55e0c861c9, 64'h17b6bdb333bca34a, 64'h000000044ea5892e, 64'h05b00c20120c8102, 64'h9ab155be32b03694);
		test(64'h75668747bf82488c, 64'h7c685eab4744ef1d, 64'h0000000770c6e286, 64'h78685c0102040818, 64'hb8b499abc44814f7);
		test(64'hef0cf60b5e140183, 64'h7cca9dc21f182940, 64'h000000000d968fa2, 64'h7008800006000140, 64'hef0cf60b5e140183);
		test(64'h58168b95ca204912, 64'h7d1e3bbc7a840d00, 64'h000000002cb3d665, 64'h1404008820800400, 64'h58168b95ca204912);
		test(64'h74172221a8e6451a, 64'hf355841804a58f10, 64'h0000000000e3838b, 64'h7050800004200d00, 64'h22217417451aa8e6);
		test(64'h105a71dfac31000e, 64'hd07f39007c34a18e, 64'h0000000006d6af07, 64'h500608000000008c, 64'ha504f74d4c3ab000);
		test(64'h26e64341334f6b4d, 64'h1c9666d7822c86db, 64'h000000001b945655, 64'h0c0620d580248219, 64'h282c76462b6d2fcc);
		test(64'hce92621b24fe0916, 64'hcac77ca70d1f7084, 64'h00000000f9606bc1, 64'h08417c8004085080, 64'hec2926b142ef9061);
		test(64'h5164efad3403ef65, 64'h1a764d46308a91fb, 64'h0000000026bd66b1, 64'h18400046300a90c9, 64'h6a7f0cc25b7f62a8);
		test(64'hbefaaea0f8409a18, 64'h336f9960808d9d2c, 64'h000000001dd530e2, 64'h3008010080840500, 64'h048f81a9afeb0aea);
		test(64'hdd04acff4b624d16, 64'hae3a3a923cdd0c0c, 64'h000000002c15c90d, 64'h0a2a02020c410408, 64'h40ddffca26b461d4);
		test(64'hb35db13fe44e3514, 64'h772a247f96556c7e, 64'h00000006d4fea94a, 64'h7720201380512028, 64'h145cb11bfc4e75ce);
		test(64'h09f23e4263e11926, 64'h43127e52996c5294, 64'h0000000003bf4711, 64'h0112604018204090, 64'he324902f9162361e);
		test(64'h368a4714b37aaf31, 64'h7f26227a7d0fb62f, 64'h0000000d8a466b71, 64'h5224025a540ba221, 64'h5ecd8cf5516c28e2);
		test(64'hc41fc6bbb9dbc283, 64'h7d76a0f2ab84b5c6, 64'h0000000223d7ed09, 64'h754680d2a0042006, 64'h13f493ee6ee783c2);
		test(64'he0e856e5231c0d2d, 64'hdd27c49a1312de77, 64'h000000030870e195, 64'h440300980000c855, 64'hb0b4c4386aa70717);
		test(64'hfa149f6eb45b860b, 64'h1fc6a551a89dd3c7, 64'h0000000345733643, 64'h15840450a8018043, 64'h5f28f9762dda61d0);
		test(64'h583f64e36580f9a0, 64'h294df6c0fce79053, 64'h000000009dad9830, 64'h214160003c868000, 64'h627ca1cff9506a10);
		test(64'h13a7af6ee1962bb3, 64'h28f3dee98ae18b24, 64'h000000002b9dd21e, 64'h28818a8108e08824, 64'h1e69b23b317afae6);
		test(64'h375d138ed2960132, 64'hb499c565e9f521b0, 64'h000000007712c4cb, 64'ha408812400212020, 64'h0132d296138e375d);
		test(64'ha87ae41ab4bea7f3, 64'h76c0b4e8f678467c, 64'h000000008746e77c, 64'h264010e8a438464c, 64'h3f7aeb4ba14ea78a);
		test(64'h427a73e6e2aaa9f0, 64'h49c7031bd1bd80a3, 64'h000000001159669c, 64'h00850109411d8000, 64'h745559f024e5ec76);
		test(64'hcb4b430b5faeb362, 64'h5b32950d99d97684, 64'h000000005c8d7934, 64'h4b32110c89186080, 64'hbcb434b0f5ea3b26);
		test(64'h0975b4b510b5e569, 64'h1f81060f0286f4e3, 64'h0000000002595bad, 64'h0281020702025441, 64'h80da7a6909ead2da);
		test(64'hf018a0d62036a1ca, 64'h25f8cbd6a9f5fe09, 64'h0000001070fa1d42, 64'h21880014a140e408, 64'h24f0e9503910c552);
		test(64'h095096e4a972b7b5, 64'h2c21cf3b554f1f9a, 64'h000000011340657c, 64'h04014238444b1b12, 64'hb1695006e5edd8a6);
		test(64'h445e0f7bdd9b2725, 64'ha8f8463bd85b782b, 64'h0000000016ffef49, 64'ha8704419880b1009, 64'h9dbb4a4ea722ed0f);
		test(64'h27eaef2b9e06a41b, 64'h7d5ebbf30336cf93, 64'h000000275dcb8e47, 64'h2952b01202220183, 64'h7f4d4e75528d9706);
		test(64'h9f3178c0bce926cc, 64'hca4f7b82ac02c781, 64'h00000000161f2f1a, 64'hc80e488028028300, 64'h6f32b4c07cd619cc);
		test(64'h85c8b268f587024e, 64'hdda1ec4b1a715fca, 64'h0000000472990427, 64'h0d816003100044c8, 64'h322592e82df51b08);
		test(64'h5ddea9cd24010ff5, 64'h0f59fcbf3ea050aa, 64'h000000037aa9b20c, 64'h044100081ea05022, 64'h0481f50f7b5737a6);
		test(64'h3e1442e517ca7a8b, 64'h549cb18839562cbe, 64'h000000001a84b3a5, 64'h109c810809520816, 64'he2ada3d45b8114bc);
		test(64'h18b79fbf67f66f67, 64'h0dd8a13a5dbcba79, 64'h0000000255f9f579, 64'h0cc0a13a18acaa19, 64'h9b9ff99b7f6f7b24);
		test(64'h337db7942bfc7d4d, 64'hdd98cab49ef376f7, 64'h00000025cd97cf25, 64'h890042349e136495, 64'hbeb2d43fed29ccbe);
		test(64'h4ef78e43be79cdda, 64'hb2bebbe58f4f08c1, 64'h00000000f7327d9e, 64'h323e1b25064d0840, 64'h8dfb4d837db6cee5);
		test(64'h7939630f7bab8690, 64'h2f37c3bc1455759d, 64'h0000000672e38458, 64'h2d35c12c10015080, 64'hf039636b0694757b);
		test(64'h55876e92e7ff1836, 64'h893625e989fc2b86, 64'h0000000013d0bfa3, 64'h881625e900c00a84, 64'h55d2b986dbff249c);
		test(64'h48ef43d44437f251, 64'h605cded64ce329f5, 64'h00000002b47d4f15, 64'h001040c64cc10141, 64'h1f2a88b3388e48fd);
		test(64'hccb86078d84232e6, 64'hea3aebc3e124cf03, 64'h00000001ae61300a, 64'h62204080c020c902, 64'h33d160e1b124c476);
		test(64'h93bd7ea2fa8f265d, 64'hdb700340e6da0f51, 64'h0000000015b9d9b7, 64'hc900034084500b41, 64'hbd51637e19aef54f);
		test(64'h85e70f580e604f0f, 64'h49d64994772cac51, 64'h000000000eda1a19, 64'h01c2400023280451, 64'h0fa44adb8f0f0d90);
		test(64'h9c1b0c3883f1c149, 64'hb49b492097b9508b, 64'h0000000016f59f65, 64'h049b002090110081, 64'h8d93c103f81c2938);
		test(64'h96c400c6d30760ea, 64'hd0d785db5a3214ab, 64'h00000000ba0cb49e, 64'hc086005940021422, 64'h0ebc756032963600);
		test(64'h4eac726c56123a42, 64'hb7dea1aed014ceb6, 64'h00000000d32738a1, 64'h8298010850108404, 64'hac8195848d39b13a);
		test(64'h399a8ff804078aab, 64'he0794d169a444f7e, 64'h0000000026780a95, 64'h0010000690040a56, 64'heaa2d0102ff2a66c);
		test(64'h9a8d767b1f4cd860, 64'h1759d32912e859d0, 64'h00000000146efaf2, 64'h1748502812005000, 64'h767b9a8dd8601f4c);
		test(64'h3c4b6b550b27fd63, 64'h42c8a76083d08a59, 64'h000000000035cc69, 64'h4040276083408809, 64'haa97873c93fe1b07);
		test(64'haa61b1099da49d0d, 64'h9a08eb8a1af73777, 64'h00000005a95aa345, 64'h0a00698202232415, 64'hb9b0b9258d905586);
		test(64'h317df0469c53e4d9, 64'h1d7d3b99d3a95550, 64'h000000027fc0506b, 64'h14381219c1091410, 64'hf046317de4d99c53);
		test(64'h80a45c0d870553fa, 64'h455a4975389ae7dd, 64'h00000000061804fc, 64'h05004900281227d4, 64'he0ca85045f3aa0b4);
		test(64'h031956e9a20d8552, 64'hfd4d6f6857328ad8, 64'h00000000159b8846, 64'h3404032801108210, 64'he956190352850da2);
		test(64'h1a8b118fa9ff59cd, 64'h5ab9d5ffca3f743e, 64'h000000f32c7d7f46, 64'h5039913fc82c701a, 64'h7365ff6af244e2a4);
		test(64'h21048902de5dc556, 64'h879d73192282eb5c, 64'h000000000882131d, 64'h8391321900024918, 64'h20984012655cd5ed);
		test(64'h7e6271ca9e02b98a, 64'h18a62d0de0539e79, 64'h0000000035990b82, 64'h08a4000140521828, 64'h4576016dc5b291bd);
		test(64'he0f6a75292b18705, 64'hada99ac5a183854b, 64'h00000000319292f1, 64'h212180c001820009, 64'hf670a45ed8940a1e);
		test(64'h069cb9b95b8ab081, 64'h1b53feeed6c1a5a0, 64'h0000000125cb1b32, 64'h024370a4c0400020, 64'h5b8ab081069cb9b9);
		test(64'h14ba271c12674eeb, 64'h7ccda280ef215ab6, 64'h000000002d181779, 64'h08418080c9211a26, 64'hb1eb84d9d83414ae);
		test(64'hc1389fe4e6f97583, 64'hc51af48eb08987a8, 64'h000000001ba75bac, 64'h050ae08690090028, 64'hf9e6837538c1e49f);
		test(64'hf3094a2242327ea7, 64'heb38139a62c9539a, 64'h000000007650d0e9, 64'h8100121062c8421a, 64'h881a06fcaddbc818);
		test(64'h7a60552a015167bd, 64'h4e70c4d139998a32, 64'h000000000dcc054e, 64'h0220804121988a22, 64'h9de70454558ada90);
		test(64'h3a0cafb9278275a6, 64'h561b8b964a7ed8cd, 64'h0000000153f082d2, 64'h10118a004074c80c, 64'hc05367f514b195ab);
		test(64'h079fd4d74e3db63c, 64'h922a857d5dabc250, 64'h000000000bd5d9b5, 64'h022801751981c200, 64'hd4d7079fb63c4e3d);
		test(64'h8a2b4fc1b60201d4, 64'h5df3345a147af0d7, 64'h000000010b31843c, 64'h0cd2000200007044, 64'hf28351d4802b6d40);
		test(64'h377f47d14118d0f6, 64'h14611a4d861e1cd7, 64'h000000000f99193e, 64'h0020024084100cc6, 64'he28becfe0b6f8218);
		test(64'hc0f049c4b353f52e, 64'h54786eca22e5d944, 64'h00000000275334f5, 64'h503048ca22444940, 64'h0c0f944c3b355fe2);
		test(64'h8895013e3312c3f6, 64'h6d4605a76458dbf1, 64'h00000000225c967e, 64'h0c06002124005bb0, 64'hc3f93321023d446a);
		test(64'hb555434f4bd4b606, 64'hbbc5be3d0b7a5eea, 64'h00000072e09fd161, 64'h8b842e2901324028, 64'h711e09e955e51f1c);
		test(64'h3ac3d320458850d7, 64'h686a4e3d466195b6, 64'h0000000039986097, 64'h4022402042001496, 64'h05d75122c708acc3);
		test(64'h5b9791416004fb1d, 64'h2c9a3b0857cf95ab, 64'h00000000b52809a5, 64'h2480000011cd80a9, 64'h02608bfd9ead2898);
		test(64'he4084bf246b00040, 64'h32e8f348eeb57040, 64'h0000000020a727c1, 64'h00c8600000100000, 64'he4084bf246b00040);
		test(64'hf65e153b697c0aa0, 64'h2159091474925ab5, 64'h0000000002e6c478, 64'h0119090000821200, 64'h500569cba2739fda);
		test(64'he16917ffd53b7340, 64'h4315d4c9a169d5a6, 64'h00000000293faed0, 64'h0211148921419000, 64'h57eccd014b69d4ff);
		test(64'h0a355cf00df0af8d, 64'hb70103969f150d92, 64'h0000000000a61b3c, 64'ha701020217140182, 64'h53f00ac5af2707f0);
		test(64'hf9f49a60d0c80309, 64'h889fb769c196714f, 64'h00000003d2acd029, 64'h0094144000024009, 64'h2f9f0659130b90c0);
		test(64'haa051904657aee6d, 64'hb437030c2f2420f1, 64'h00000000030ab5ad, 64'h2435010c0e042061, 64'hdd9e9ab52608550a);
		test(64'h0334df3d938c74f0, 64'h0ecfc1c6251a5019, 64'h000000000113915c, 64'h068300c4201a4000, 64'h3eef3803f0b84c63);
		test(64'h21c5a0e1203542f9, 64'hfb2eb91b2b02b63c, 64'h000000008960601e, 64'h4800310900023624, 64'h9f2453021e0a5c12);
		test(64'ha3d2d1bef39ebc50, 64'h73b3b96b940c9528, 64'h000000002ed576f8, 64'h70b0b84b80041000, 64'h9ef350bcd2a3bed1);
		test(64'he86c53345ea0c602, 64'hf86dc08908f0470e, 64'h00000000077c8d71, 64'hd040408000c00004, 64'h392b1cc50ab58093);
		test(64'h705444776611a400, 64'hc2e36d8d36a48748, 64'h0000000012247630, 64'h80c0208904000000, 64'h54707744116600a4);
		test(64'h739244cd2d8d1c46, 64'hd601188dd8e5d7fe, 64'h00000001a3c66623, 64'h4200180c1840d08c, 64'h91347278731186cd);
		test(64'hf156036a077c23d1, 64'h5b5c250297ac0fd6, 64'h00000000674cee7c, 64'h0154250201040e82, 64'hc0a94f95c847d03d);
		test(64'hc0727fec3ce86249, 64'h41934201d35a00cd, 64'h00000000004d894d, 64'h4110000181080041, 64'h1b0ccdfb4dc36819);
		test(64'h94b45250097d278c, 64'h41710a762f51bec3, 64'h000000000cd13d38, 64'h002008760901b0c0, 64'h92d2a4a009eb4e13);
		test(64'h00f9f172ba44cd7e, 64'h2c46a62fe164db64, 64'h000000000992abaf, 64'h0c420404c0609b60, 64'hab44dce7009f1f27);
		test(64'h401ca54feb584bd2, 64'hb0356558346c4fc5, 64'h00000000033d95bc, 64'h9014450010244d04, 64'h08c2a5f87d4a781e);
		test(64'ha28372cd9adbc61a, 64'h2568ebaca1f0b716, 64'h0000000081ab9b35, 64'h2060a98ca0300304, 64'h8d738ac293a4a6e7);
		test(64'hb2b66195358c53f8, 64'he32c23b39c32b55f, 64'h00000002d6d54178, 64'h4124030304103558, 64'ha9866d4d1fca31ac);
		test(64'haebfa68d6ee667f5, 64'hf454d5feeda8f67a, 64'h000000ab9467b37c, 64'h844451dc6180f652, 64'hf59db99b27a9efab);
		test(64'hd280175996ad7916, 64'h3645b03e6d34a664, 64'h0000000014160aa1, 64'h124120346c100460, 64'h69da97612d087195);
		test(64'h73856974645bd628, 64'hbb7f737337abeb84, 64'h000000d85cf287c8, 64'h9a462052368a2200, 64'h3758964746b56d82);
		test(64'h3ae1bb30fce8dd53, 64'h5a55d2fcccde3829, 64'h00000001e6ccfd19, 64'h0a5512a0c4ca1009, 64'hd4fca3eed2353077);
		test(64'h5e29d46899feae19, 64'h79de4b9208aff505, 64'h0000000161207ea9, 64'h218e4b82008e1401, 64'hda618e4966dfd562);
		test(64'h14e8a1546ebd4baf, 64'h51762854b5b73af8, 64'h00000000b1757a75, 64'h01560814a4853278, 64'haf4bbd6e54a1e814);
		test(64'h1a6b6b044357ea8d, 64'h9eb5325cef4a4618, 64'h000000006a68a3b5, 64'h1031105cca400608, 64'h046b6b1a8dea5743);
		test(64'h9d5acb6665ee5494, 64'h12165b9042582d3d, 64'h0000000002b72a4a, 64'h02161a1002100828, 64'h868adda9997c5ae6);
		test(64'hee2f799c153e7227, 64'h84859b5562ca6703, 64'h000000000db581eb, 64'h04041b4160402103, 64'h774fe9938ac7e44e);
		test(64'he544858e906c530d, 64'h0f46855fcdefe8eb, 64'h0000001773a0f105, 64'h034201018c24c029, 64'h63900bac227a171a);
		test(64'h92654f3d2f676dfa, 64'he5fd2dbf5a1f9da1, 64'h00000083377a673e, 64'h25a42d334a0d9d20, 64'h1f9b9ef5619a8f3e);
		test(64'he628f280854ceada, 64'hde5287a24139858f, 64'h000000003315129a, 64'h0a1006224028848a, 64'h1467014f32a15b57);
		test(64'h8b8f74cc91e37544, 64'hf3a6f657dbe962ae, 64'h0000008edea53dc2, 64'hc304425453a12008, 64'hcb46115df2e2331d);
		test(64'h875791971585dbeb, 64'h060c7a8b749d4a9c, 64'h000000001a4b39fa, 64'h04086009648d488c, 64'h79197578bebd5851);
		test(64'hd42e76da42675709, 64'hb317df4572197be7, 64'h00000028cda49ac1, 64'h3102094070113821, 64'h42e6ea902b746e5b);
		test(64'h57a62c5af07f50d0, 64'hc26a481284b39a71, 64'h0000000001abcf4a, 64'h006a481080809200, 64'ha0e0f0bf1ca5ab59);
		test(64'h1b1534917c184105, 64'h96b4b485715e90c7, 64'h0000000029bde605, 64'h9680140020040005, 64'hd8a82c893e1882a0);
		test(64'ha513ae9a064cfc26, 64'h0e7f12786647ac5e, 64'h0000000089a679e3, 64'h000c10302646040c, 64'ha6bac45a983f3190);
		test(64'h10f39b5a1be7f486, 64'hb072b8ed1d63daef, 64'h00000007ed4dfe46, 64'ha04030ec0d634206, 64'he7d8612fcf085ad9);
		test(64'h6c4e0c9369c6469a, 64'h1e5635c6af792c97, 64'h00000003594b303a, 64'h0c520580a2182092, 64'h30c9367262599663);
		test(64'ha28c8e15efe21b0e, 64'h6c34503bc6aadcb8, 64'h000000002113fa61, 64'h6434502100a280b0, 64'h0e1be2ef158e8ca2);
		test(64'h7a81ceb00e05a701, 64'h820dd7cec38e4c0f, 64'h0000000027681111, 64'h00058046408c0001, 64'h815e0d73a07080e5);
		test(64'hf7c50f9712b5b357, 64'h52afcd37fc74edf1, 64'h000000f29de23d2b, 64'h408e0825ac3064b1, 64'h73ab217a0f6bfbca);
		test(64'hebe706cea3dd586a, 64'h55086a931275b85a, 64'h00000000090d373b, 64'h05084a8210603048, 64'h3b09bdbe9a5277ac);
		test(64'h217280a4156005aa, 64'hed9cc5f1dbbcef21, 64'h0000001291425016, 64'h440084b00008ca20, 64'h2a900a5512b14058);
		test(64'h033e2ed3b7aa7ebf, 64'he644fb8c7e896582, 64'h000000000a5a37bb, 64'ha444d2807e086582, 64'h0ccb8b7cedaadbef);
		test(64'h44accf8f470f57c9, 64'he6a77c7b46e19b26, 64'h000000057263f158, 64'he481603a42619102, 64'hd1f0d563113af3f2);
		test(64'h80263252984e5190, 64'h35d37028b6bea933, 64'h0000000002650714, 64'h10c02008a2228100, 64'ha8909127c4a41046);
		test(64'hcf04f08d6c1df8a1, 64'hbedeeaeb588fcb10, 64'h0000001385c96b78, 64'h34cc02cb58028010, 64'hf08dcf04f8a16c1d);
		test(64'h6eb62fa575a21086, 64'ha2322fa87f93b527, 64'h00000001ffeeb446, 64'h20320b2010802006, 64'hae450861766df4a5);
		test(64'hba3dd450ca3f3b8d, 64'h45aca4a50e6006ba, 64'h00000000003d0ab2, 64'h402ca4050a600032, 64'h27cecf3a5071c7ea);
		test(64'h3a5dcc378cc42837, 64'h95742476cc9f4da7, 64'h000000012d7dc88f, 64'h9414006080140187, 64'h312314ec5cba33ec);
		test(64'h01e4d6dd1a99fafc, 64'h8cc3787ed59ff609, 64'h00000001957139f6, 64'h88806826159af600, 64'hd802eee96625fcf5);
		test(64'h951a599866426ba5, 64'hd060113bc704a632, 64'h00000000014d8e2c, 64'h1000002343042022, 64'h9ea599185662654a);
		test(64'h1df22dc2229963fe, 64'ha27ea4b4f1896eb9, 64'h0000000072e09f3e, 64'h8022203051006eb8, 64'hfd936611c11ef12e);
		test(64'ha3e4453d33aef224, 64'he2099ced31b1a6c0, 64'h000000001609ff34, 64'h820914cd20808200, 64'ha3e4453d33aef224);
		test(64'hf56a74685879758d, 64'hd9a3c1d330694426, 64'h000000000eb243fa, 64'h80a3015220600422, 64'h256d5d725fa91d29);
		test(64'h89f9dd291a805f2e, 64'h3c33810b4b675410, 64'h0000000000b7ac0e, 64'h280000024b425400, 64'hdd2989f95f2e1a80);
		test(64'hd7e410fa53d69eb8, 64'h0d3bae36ba0b9d85, 64'h00000000e00d2af4, 64'h0111aa148a0a8d00, 64'hbe8d025f3a9ed647);
		test(64'h7f06cfd5b1d44bfe, 64'ha5884ca95f08dce9, 64'h000000001cf2895e, 64'ha00848880900dce8, 64'he872fd8709bfeacf);
		test(64'h1648f5bf7a3cd710, 64'hc174c6f3c4636abe, 64'h00000000475e9248, 64'hc074407244216020, 64'h04d73cadfe5f2194);
		test(64'h8f1f47ced1b0c3eb, 64'hc6af207f490638ac, 64'h000000002cf4ea0e, 64'h402b000c0106308c, 64'h0b1dbe3cf1f8ec74);
		test(64'h337fead20eb59fdd, 64'h0f1c883bf370a3a2, 64'h000000000fea09dc, 64'h0314082993708382, 64'h0be56f77ccdfba78);
		test(64'h1c55582c9800ea65, 64'h634bd23779a4d2f1, 64'h0000000025a861ad, 64'h020a000038841221, 64'hd59a6400a41c2caa);
		test(64'h57ccef03ea150714, 64'h5d735ba11856681a, 64'h00000000370b9584, 64'h4901120008502010, 64'h0cbf335d410d45ba);
		test(64'hdade73a5866b824a, 64'h395fd973285287ce, 64'h00000001be6a4b4d, 64'h1806513200020244, 64'hb7a75acde992a182);
		test(64'h7df64bb5a8d81141, 64'h4b4e101855e3d123, 64'h0000000006da0c19, 64'h0146000001028001, 64'h51b18828ebf62dda);
		test(64'h897d4fa11b1a3e41, 64'hdcffceccac91ba7d, 64'h00000093ebe093e1, 64'h902348488091a201, 64'h28d3527225f8eb64);
		test(64'h0abc5a3b6a7ba649, 64'h02cd2c053005e345, 64'h00000000006c99b5, 64'h02c9280410044101, 64'h50c75a73597b9568);
		test(64'h84201ffab4f399c3, 64'h693ceb7ed2246e30, 64'h00000000103fb510, 64'h21286a38c0244030, 64'h99c3b4f31ffa8420);
		test(64'hdb0bc1e37e85aaec, 64'h20ae99f0993d9ab9, 64'h000000001679877a, 64'h00ae881018291a30, 64'hdc554abdd3c207e7);
		test(64'ha5f2a3be5ba66fcc, 64'h345064fda3555013, 64'h000000000babc650, 64'h2450206523541010, 64'h5cd75af46f33ad56);
		test(64'ha6d201bd1ba39e73, 64'h34319cf6b1a3258f, 64'h00000000a82e3f43, 64'h0030988681a20583, 64'h4b65bd80c5d8ce79);
		test(64'h2f0eb52690b0e004, 64'h9fa4e8acec2100c4, 64'h0000000001e69611, 64'h0580288000000080, 64'hf2e05b62090b0e40);
		test(64'h2d312c817a2bf3c5, 64'h8b375974669ff562, 64'h00000005c90697ec, 64'h011710242699e042, 64'hda8efc3587c48324);
		test(64'hacc0480b7313d208, 64'hecc112a5341877ac, 64'h0000000017c0eaa2, 64'h8c00102524004080, 64'h3137802d0ccab084);
		test(64'hf194727e2e1e2c43, 64'h7e81205051f760db, 64'h000000001c5c0e53, 64'h3800205040542003, 64'he7e492f82c438747);
		test(64'h224afd15d123d8da, 64'h526c05661abae9eb, 64'h0000000035944eb6, 64'h504004200aaa0962, 64'h4cb8b5b125448afb);
		test(64'h5c1f0dac28f886f8, 64'h0795610dcdbdc9f5, 64'h0000000239c4f23c, 64'h0011000dc08189e0, 64'h944f414fe0c5caf2);
		test(64'hc8f5b1dfde266f26, 64'hd32d9d4571152a78, 64'h0000000062f3e974, 64'h9320850151140830, 64'h266f26dedfb1f5c8);
		test(64'h12460ee427aa9e2c, 64'hac37120ad6a7c010, 64'h00000000000c83d4, 64'ha8250200d4058000, 64'h0ee412469e2c27aa);
		test(64'h067581be85d88b90, 64'h1c61eaa0228dde87, 64'h0000000007c33258, 64'h0421a8002004d200, 64'h60ae817da11bd109);
		test(64'h2b2f71f3739b84fa, 64'hbfe53bba99e4cd73, 64'h000000567cf5625e, 64'hb9a50b1898040d62, 64'h12f5ec9de8fc4d4f);
		test(64'h800d54c37c183829, 64'h08ade6e0bfd92219, 64'h000000000eacf0d3, 64'h08ac02800e010201, 64'hc3a80e40163424bc);
		test(64'h90ea4ba3c097361d, 64'hc78187e63a7a3f31, 64'h0000000211d40bb3, 64'hc6000122306a0321, 64'h392ec06b875360d5);
		test(64'h82c3e4e66179270f, 64'hd29238bf3a11f681, 64'h000000004d99a32d, 64'hc00218a422110681, 64'h41c3d8d992b61b0f);
		test(64'h3c2b29d25490552c, 64'hdaaefc95a385be86, 64'h0000000334ac0852, 64'h108a240021048a80, 64'h3ce8688715065538);
		test(64'h65df8c8f768bd47b, 64'h68539ea3ca3abd13, 64'h00000001bed6a757, 64'h48518821c8281d03, 64'h131f6abfb2ede61d);
		test(64'hcbe6416c8df1eca9, 64'h8d2a6d7b1f640530, 64'h0000000036c746ea, 64'h050a683a19200410, 64'heca98df1416ccbe6);
		test(64'hc8116571b289813a, 64'hbe7baad1fadb9cb8, 64'h00000090947b6587, 64'h3833088098010c90, 64'h3a8189b2716511c8);
		test(64'h67f4ee1d975c0581, 64'h9f5cc5c80057fdca, 64'h000000003ef1e038, 64'h925885800000b002, 64'hf19d47bb536d2405);
		test(64'h1b78fa6bbb7360b1, 64'hc8025f88c8ab8a30, 64'h00000000005d3563, 64'h8802468800098010, 64'h60b1bb73fa6b1b78);
		test(64'hc2d5a52c20d65124, 64'hf475cf3aee2b3486, 64'h0000000c5e5a2092, 64'hc0200d1848082080, 64'h83575a3808974518);
		test(64'h22bd588f7174836f, 64'h5726aa7a018951a9, 64'h0000000001621c17, 64'h02262040008850a9, 64'hb8b29f437e114fa4);
		test(64'hf0524249af7f094a, 64'h3bf944dcc97ae5d8, 64'h0000000c292afe15, 64'h235940dcc010a090, 64'h494252f04a097faf);
		test(64'h23d4fd9cbecc6613, 64'hf43cd4458c541a1f, 64'h0000000008bebd33, 64'hf418500180500013, 64'h39bf2bc4c866337d);
		test(64'h74602f173adfd5eb, 64'head97e18b8e27080, 64'h000000001885e7db, 64'he2517e0828e05080, 64'h74602f173adfd5eb);
		test(64'h7f3da3e9d7dd9461, 64'hfa969b166f891709, 64'h00000000fb4c4ff1, 64'he8968b060a011001, 64'h3ebfd653eeeb9268);
		test(64'h5532b9af4d3ce767, 64'hbf52de4f8ea1a769, 64'h000000055d8f65fd, 64'h3d02924c8c218629, 64'h3c8e9bdb31aa5f76);
		test(64'hd6db03b4b1f61e67, 64'h2a82031c71e88b9b, 64'h0000000001fafcc3, 64'h0282030c00e8030b, 64'hd20cbdb66e87f6d8);
		test(64'hf6420a8e9ac2dc4c, 64'h4ab727f6f921caf4, 64'h0000000a114731c9, 64'h4a23058269200860, 64'hcdc4a92ca0e86f24);
		test(64'h7953a0dc0d3db461, 64'h6f2028b4a254f749, 64'h000000001cab0ee5, 64'h2a0028a482441401, 64'ha3b6ec503e0e9278);
		test(64'hc9ed500e990aace7, 64'hd7787c3753f3607e, 64'h00000031da194273, 64'h1648480242b0604e, 64'hdb3aa066b0057b63);
		test(64'h0f8430631fff593e, 64'h0eecd9599d29280c, 64'h000000001e2497f7, 64'h0eecd91184092808, 64'h48f03603fff1e395);
		test(64'h5ebee798b3e0f95c, 64'h5747a122baceefae, 64'h0000000f373b8f26, 64'h41062122804e8aa8, 64'h0bce356fbeb526db);
		test(64'hc10a127d221759f1, 64'hf8e45025e0bf2b02, 64'h00000000180792ea, 64'h10041024a08f2002, 64'h340a48d7884d56f4);
		test(64'h29d1ee43ca7cd5d4, 64'h5c7534edfa99d97f, 64'h0000002ad4736ed4, 64'h101520a1f0914954, 64'h2bab3e53c2778b94);
		test(64'h4e4e22c3162f550d, 64'h520f8e6920b9e8e7, 64'h000000005e192d05, 64'h0206046900914025, 64'h68f4aab0727244c3);
		test(64'hfcd0ec16647242f6, 64'he922bc30ab92dbf3, 64'h00000003c6d434be, 64'h89008430088013d2, 64'h24f662e47386f3b0);
		test(64'h7ff90a0ab0056284, 64'h07613c689aef4941, 64'h000000001f91c0b0, 64'h0400004818240100, 64'hbff60505700a9148);
		test(64'hce7bc52ad606e793, 64'hf2189f1703d96e9c, 64'h000000019e5281bc, 64'h620880060389620c, 64'ha25cb7ec397e606d);
		test(64'hf71c673f00d4fb41, 64'h9b5bd92c916da2f7, 64'h0000000db13c4ba1, 64'h9a001824016ca081, 64'hdf82002be6fcef38);
		test(64'h8e90f9656f9d2472, 64'hc8e0e13563f142ba, 64'h000000002cfbf98d, 64'h88e0813102404288, 64'hd881679f95f6602b);
		test(64'h56cc7bb3404f4ebf, 64'h1732de0ae30f9fe2, 64'h0000000383aa3ceb, 64'h15000402e1038be2, 64'h101f1bef5933deec);
		test(64'h86b5e8cbb668385d, 64'hb5aebf3802db5f6d, 64'h00000025ad06a317, 64'h11a63310000b0269, 64'h4997ea43a7947c4d);
		test(64'h3ab673d48ac29293, 64'h03b6f90a67cdd376, 64'h00000005f74162c5, 64'h0220a90005089046, 64'h86c6a283cd17ac9e);
		test(64'he81eeea890b85550, 64'he32da10a06d271fa, 64'h0000000038da2ad4, 64'h4009a00002422140, 64'h5055e260a2bb4bb2);
		test(64'ha78528ea3f4eeb99, 64'hbd26942e85e5b00e, 64'h0000000033435ab4, 64'hbd04142681643002, 64'h52daab28b1fc66eb);
		test(64'h6b4a2d1c665fb8ee, 64'hcb9c0e55c65efc1f, 64'h000000079667fdce, 64'hc0900c11c64e1c0e, 64'h38b452d6771dfa66);
		test(64'h7d24502e69a0a627, 64'h4a8f4d1d54c88eab, 64'h000000006243496b, 64'h488308011048020b, 64'h50694e5642eb47a0);
		test(64'hdefc2564e77bd576, 64'h6b150d25f456bf5c, 64'h00000002d9eeed5d, 64'h0b010c25b4449718, 64'h4652cfed675db77e);
		test(64'h6ab42b3cf7be4522, 64'hcb4d4068cb343128, 64'h0000000001c47be6, 64'hc94d002009040020, 64'hbef72245b46a3c2b);
		test(64'hd0fe7aaa771f134a, 64'hdbd66e987984bfec, 64'h00000038ff6f526a, 64'h9254681870041a48, 64'hf177a431ef0daaa7);
		test(64'hc0fe14202483cd93, 64'hcb5c9f86a01bcec8, 64'h00000000c7a813f4, 64'h0844018600198448, 64'hfec02014832493cd);
		test(64'h7e38b7f044db4b55, 64'h0c3cc5c0eaec8883, 64'h0000000007d7a349, 64'h0818c18088c88081, 64'he7c1def022bd2daa);
		test(64'h37f5533a63af1152, 64'hea4b067da9665bf0, 64'h00000000b2b8ae95, 64'h8a01062d80404920, 64'h115263af533a37f5);
		test(64'hfffe3b8f16526b47, 64'hb51165ee2d2efe51, 64'h00000007e59c85ad, 64'hb00124482124d051, 64'h374ffffd978b29a1);
		test(64'h6a8933094adb17ed, 64'hd8bcd28b7972fa82, 64'h00000001646b2b16, 64'h481450894132ea02, 64'h9a26cc061a7e4db7);
		test(64'h8fd4be039380fff7, 64'hd3f23326acf6e3c8, 64'h00000004f5c620fe, 64'h524230000cf6e2c8, 64'hd48f03be8093f7ff);
		test(64'h0257cba8f870fc0f, 64'hd8cbc5725650fe37, 64'h000000002f533fc7, 64'h08ca01600650c017, 64'h3ff01f0ed31540ea);
		test(64'h286b36ad5d13320b, 64'h8e49aa7cc87af6af, 64'h00000004eab6534b, 64'h8a08a844084a200b, 64'hc8bad04cd614b56c);
		test(64'hc45adc11e0864882, 64'h3d65064b62e32493, 64'h000000000288748a, 64'h0040024102020002, 64'hb38832a521147016);
		test(64'hf91162386449a61a, 64'h5024a63bd587f3d6, 64'h000000018bc50d45, 64'h002404088504c0c4, 64'h892c6f449aa41961);
		test(64'hf30e6067aec8c9b1, 64'h1e5705b7e2551462, 64'h0000000024c2f702, 64'h1646010640511002, 64'hab3236e4fc0b909d);
		test(64'h8b014ebf77cce6ca, 64'hb99fc0817dcd8d87, 64'h0000000260bf7eaa, 64'ha98f80014d0c8882, 64'hd18072fdee336753);
		test(64'ha0c18b2d935d975c, 64'h72ee2ade5b117b72, 64'h00000004c18cbcba, 64'h6288289c51016960, 64'h6d536c572e87a034);
		test(64'ha2249350869fc504, 64'h0d26ef020fdf3b8e, 64'h000000006866be12, 64'h010064020fc22008, 64'h188a05c6f6921053);
		test(64'h962f155b578da679, 64'h9ac61a5db06e0375, 64'h0000000069ce935d, 64'h88c6005520280361, 64'h956bbae4a27a96f1);
		test(64'h372f16c99486a233, 64'h447e2c93752f43b7, 64'h000000015cc98c9b, 64'h044a0400642100a3, 64'h45cc29616893ecf4);
		test(64'hb58a7a74d18310f0, 64'h28391c706f582ad1, 64'h0000000008b7840e, 64'h0018003004082a00, 64'hb5b87a4520f0e243);
		test(64'hf4d0c614415e0ec4, 64'h388d95acf83583d9, 64'h00000000d1428658, 64'h100084ac00348210, 64'h28c9e0f8c80dad82);
		test(64'h7e52430361e23e9e, 64'ha09cfb9a62bb9d63, 64'h0000000288c764e2, 64'h208c0b80403b1162, 64'h6874c797e7a42c0c);
		test(64'heed57ec92e07d299, 64'hc6f1cc4771045b7c, 64'h00000000fdbca746, 64'h04e0004750004864, 64'h992d70e29ce75dee);
		test(64'h5ec1bb1d2c0b0cca, 64'hdc33b0b3a5af6853, 64'h00000001e3cac59a, 64'h4412001180294042, 64'hdd8ba7380335430d);
		test(64'hb46d07e6c0b24243, 64'hec262f98c5e5d607, 64'h000000015c79944b, 64'h60000b0804044003, 64'h2db6e067034d42c2);
		test(64'h1312f2fccf0d7c6b, 64'hae41454962e71c53, 64'h000000000126a2fb, 64'h2e00014122e01843, 64'hf4f38c84e36d3f0b);
		test(64'hf46aed18e739a6ab, 64'h6ca23a8a12071f26, 64'h0000000006ba4935, 64'h6822228200061506, 64'hdb6c9aea1fa97b24);
		test(64'h17d2563b55301898, 64'h7067cffad1dd5ea9, 64'h000000192c7b90ca, 64'h30468a9800181280, 64'h30aa6424e12b37a9);
		test(64'hc15e551224546e54, 64'hd89cd8203fddd388, 64'h00000000c7648d28, 64'h1010480023589100, 64'h5ec112555424546e);
		test(64'h9fd78b2b26f98a2f, 64'h7a38750dda6512fb, 64'h00000000e8343a97, 64'h6208550c5021005b, 64'h4f15f9464d1dbe9f);
		test(64'h8fcb0849f6f6061e, 64'h8aeb8249437dad92, 64'h000000007dcfba13, 64'h8a638209000c0590, 64'h02162f3e094bf9f9);
		test(64'h25b299365fb07249, 64'h82b2d8d09080a0ed, 64'h00000000003ecb55, 64'h80a008c010002021, 64'h07fa681b17a19366);
		test(64'heeb1907d704c3aec, 64'h59177ff72dcd9999, 64'h00000054907b0e6a, 64'h5912704601c49890, 64'hbe6072dddc358cb0);
		test(64'h25704efc8a1744ea, 64'h2cf4bc9f3f8910e3, 64'h00000002b87e145e, 64'h0410808e22091042, 64'h158e22754ae027f3);
		test(64'h91a0168475aa5a02, 64'h6054c02ec0fbce36, 64'h000000000009acd1, 64'h4044802480590004, 64'ha5805daa9412460a);
		test(64'h8da20e9f321b742a, 64'hdbf2c343f4a30842, 64'h0000000025a93319, 64'hc212424340210040, 64'h27a80b6fc84ed18a);
		test(64'h93c5fdac07241ed2, 64'h174cb65d5129a26f, 64'h00000000bbe31862, 64'h000c841001292222, 64'h24e04b78a3c935bf);
		test(64'ha405391d80788aeb, 64'h8b21ac0ff67ba13e, 64'h0000000216d83c95, 64'h0a0000078412a116, 64'heba22d02746c501a);
		test(64'h9b1714d4b0a0d9fc, 64'h4af4cc55e456674f, 64'h000000018c7a823c, 64'h026008402414274c, 64'he8d92b28050d3f9b);
		test(64'hcaa5a1e3666cf841, 64'h830db798877411f1, 64'h0000000033c636c9, 64'h800c330887001001, 64'hf482999c52d3c55a);
		test(64'h81e488b9a264a592, 64'ha7cbe2fa4c094859, 64'h0000000047117004, 64'h2083205044080808, 64'h7644d842615a9851);
		test(64'hde78a5bd4ada6c89, 64'heea504747f65da10, 64'h00000000dd2f2a14, 64'h448500641b041010, 64'ha5bdde786c894ada);
		test(64'hf7a837d0dee795a4, 64'he018e0435315b38f, 64'h000000000e99ceb4, 64'he008c00350113104, 64'h15ef0bece77b25a9);
		test(64'hab83e66890fe9b28, 64'h05df33a6f520ac1e, 64'h0000000061d249a4, 64'h044133a231200810, 64'h299bc2ea28e6bf06);
		test(64'h97dd701cb0ee2ac6, 64'h8e37b576797b8713, 64'h00000016d6199b12, 64'h8c13016641298012, 64'he0839ebb4536d077);
		test(64'he9333fb81230d4dd, 64'he4d25cf1b0d22234, 64'h000000001c6f6243, 64'h8402406120502224, 64'h4ddd2103f38b9e33);
		test(64'h4a6eb4c5359d8b70, 64'h616b2da6b1366c66, 64'h000000009eaa762c, 64'h014921a280262c00, 64'h5c76e20da1b91e53);
		test(64'h8c38bcf0ce3fd93e, 64'h4a6b5e99096a290c, 64'h0000000004c764ef, 64'h4a035e8900422908, 64'h83c80fcbf3ece39d);
		test(64'h3f6d46ed586f3e5e, 64'h8ee9718c119fb7a2, 64'h00000000ef8f1ef1, 64'h84c0308c101f13a0, 64'h529fcb5bcf9719b7);
		test(64'h25287312d83f204d, 64'h539690d8ccd4ed4d, 64'h00000000104b8c8f, 64'h518000d8c0800849, 64'h41a1123bf34ee801);
		test(64'ha42f39efba71b7d7, 64'h95ed74184d624178, 64'h00000000147b299a, 64'h912c140845620138, 64'hd7b771baef392fa4);
		test(64'h79867bc0dab3dbfa, 64'h8f3c8549891502cd, 64'h000000000244cd7c, 64'h0a308541811502c4, 64'h946b0c7b375e5f7e);
		test(64'h21ad613f880e3b88, 64'h86ade2ddb81fc5ff, 64'h0000000fb1f2e188, 64'h06ad020038038588, 64'h11dc7011fc86b584);
		test(64'h48684137374965b4, 64'h35ed750193361a7f, 64'h000000001c8dc034, 64'h30cd210011220a34, 64'h2da692ecec821612);
		test(64'h21a8e05b8dcf098b, 64'h905b868e82979558, 64'h0000000000916b89, 64'h901a068800830118, 64'h5be0a8218b09cf8d);
		test(64'h65a8d3c81038ec72, 64'h9bf7553711f9c12a, 64'h00000000686823b5, 64'h0040150310c1c008, 64'hc240d8b3a295327c);
		test(64'h597f677849df3828, 64'h29c51d9031378c58, 64'h0000000003734bd1, 64'h01c11d0031008400, 64'h78677f592838df49);
		test(64'h6060affa47bdf540, 64'hc4f31d0c5fb3deaa, 64'h00000004c3d3f7a0, 64'h84201d045bb14800, 64'he71d10f59090faaf);
		test(64'hc1b3938b77005397, 64'h43862f81066856f0, 64'h0000000002d1f8d9, 64'h4200008004284270, 64'h53977700938bc1b3);
		test(64'h41dfca0ce0153a5d, 64'h6cabdd0215022769, 64'h0000000008be80ab, 64'h0002910211000561, 64'h2ad0ae35ef820cc5);
		test(64'h061fa204a782d967, 64'he289a237df7d6515, 64'h00000000be48e04b, 64'h8208223016646015, 64'h158090f26eb9b514);
		test(64'h59b5411b36067a9f, 64'he75d96da2df331aa, 64'h00000008ac0f416b, 64'hc619800a05d101aa, 64'h09c96fdae5564e14);
		test(64'he8a8d86179c3fd49, 64'h8f2cd67ba58008f3, 64'h00000000637315d1, 64'h8e0c807ba1000821, 64'hfb29e93cb1687151);
		test(64'hded402209b935422, 64'h3ccd989a20e13a0a, 64'h0000000003e80251, 64'h1c08908820002008, 64'h717b80086c6e8851);
		test(64'h4cbf76617e533afe, 64'hdd0721658928e30b, 64'h0000000005bda836, 64'hd10201418820e30a, 64'hdf2368e6ace7f7c5);
		test(64'hb799efa63479100d, 64'h6d8f7bd3c68e416d, 64'h00000005e7791207, 64'h280d0b8204000029, 64'h6b83e00266b795fd);
		test(64'h51f8fc7947e0a6af, 64'h38b3880a01d72c22, 64'h00000000005cee17, 64'h3800800800c50c22, 64'h1db0a9af54f2f3d6);
		test(64'h1260a697106fcafa, 64'h469899d60b3cebef, 64'h0000000111717b7a, 64'h460080140b3849ea, 64'hf6085f530648e965);
		test(64'h6d08f6dbe69d89f8, 64'h290ca307dedbcceb, 64'h00000003dcf3b6bc, 64'h290c03025a824ce0, 64'h9b76f119016bbdf6);
		test(64'hbcccbc7d5d6c21b2, 64'h08eb602ed20ad571, 64'h000000000e8f3416, 64'h08a320204000c510, 64'h1271ae9c7cbe7ccc);
		test(64'haa11c8702e83bc9b, 64'h764fc17ee3e6fd22, 64'h000000121dc1a379, 64'h6002c12062e44c22, 64'h8b2ce36eaa4432d0);
		test(64'h350cad4c488a3858, 64'h7dcf0529c1ce3a28, 64'h0000000036669579, 64'h48410100c1021800, 64'h8a4858380c354cad);
		test(64'h4e84a4667e3e2c5c, 64'h2d518af376cac704, 64'h00000000308d7cc9, 64'h2d5002f026024600, 64'he4484a66e7e3c2c5);
		test(64'hebf30f0e5d62138a, 64'h49505771b177752d, 64'h00000001f381e454, 64'h0110526020116024, 64'h19ea54323f7dd0f0);
		test(64'h7802df4700637087, 64'hf5c61a6b17e377a6, 64'h0000000e0f983f8b, 64'h3400002806e01026, 64'h00c90dd22d80f7d1);
		test(64'hea2ac1ad667798c9, 64'h1409f731993465b8, 64'h0000000005868709, 64'h0009353109006088, 64'hc9987766adc12aea);
		test(64'h1d846ccffd4e6373, 64'hc1bc52c47ba84375, 64'h0000000018cfe9fd, 64'hc1a840c418280345, 64'h393befd8c9fce284);
		test(64'h63673648cc476eb3, 64'h639a303bf88e2cae, 64'h00000000f1c993f9, 64'h60901003b08c2486, 64'hd133ceb9d9c9219c);
		test(64'hcebea777df8fdb77, 64'he21aad6edaaaf901, 64'h00000001bf7bfdef, 64'he01aa82eca28e901, 64'hcd7d5bbbef4fe7bb);
		test(64'h8777fdd46be7ccb3, 64'hacaf6ce35c814fea, 64'h00000004aff8af95, 64'h80a56c235081058a, 64'hbd9eec33dd2d71f7);
		test(64'h834a46507c7cf7f5, 64'h588ff3c2fbf3535a, 64'h00000002924f1cfc, 64'h1001f042e3d35312, 64'h50191a2cf5fdd3d3);
		test(64'h20719293ae43237c, 64'h532d5be489ccfa3a, 64'h000000002551909e, 64'h522542048080da30, 64'hd38c1cab6c68d480);
		test(64'h2b303005f63aad4e, 64'hf2d4a277b1fc4b94, 64'h00000001490bc729, 64'hb2c4803521684190, 64'h0350b203dae46fa3);
		test(64'ha796311f04f9d603, 64'h1530c6a8b49bc56f, 64'h000000003408f783, 64'h001006a814898003, 64'h9f20c06b69e5f88c);
		test(64'h3ac96cc729e44925, 64'h42af85ea866f68f7, 64'h000000034ac8d295, 64'h428501e080222045, 64'h92a4942736e35c93);
		test(64'h526cbbc3f26b6be6, 64'h1c95e8568b4b84b1, 64'h0000000010ae6bcc, 64'h1081a052824b8030, 64'h97d9f19777c3a19c);
		test(64'hae470f19bbda1ff8, 64'haf1f0bb8965b55c7, 64'h0000000f8fcf7cf8, 64'h861d0b30801b55c0, 64'h75e2f098dd5bf81f);
		test(64'hdc76ff75fe4272ac, 64'he3e6e6d371e5dd49, 64'h00000030ffb790c2, 64'hc2e6e08041c14940, 64'hb9ecbaff81fd5cb1);
		test(64'hdcbeda4edcbe64b3, 64'hd84dabca0b7c54ba, 64'h00000001ed678fbd, 64'h504c23c80310448a, 64'hec91eb731b7aeb73);
		test(64'h6b0f16a14fcec293, 64'h9a84c441111f9bd6, 64'h00000000034aba55, 64'h9a84044101108886, 64'h944ae9f083c6f1b3);
		test(64'hfd54b0ed05639161, 64'h6f5c6923a9a72e03, 64'h00000000f7528ac1, 64'h0114402308052001, 64'hfba2d07b0a6c9868);
		test(64'h3be229d063c1809f, 64'h55e393088bc9c45e, 64'h0000000017c23d8f, 64'h40e200088000805e, 64'h07688becf60243c9);
		test(64'h2927273c50888056, 64'h94b5187193af44d6, 64'h00000000058c940f, 64'h8401002010004094, 64'hd83c68d802950522);
		test(64'h8f74bbd7ac7defdf, 64'hbdb7118ea62503c0, 64'h0000000013b9df7f, 64'h30b6118aa62103c0, 64'h8f74bbd7ac7defdf);
		test(64'hceb8ec63e1dfb9c7, 64'h2063b4ed88229774, 64'h00000000026b3399, 64'h000394e988009434, 64'h9b7c1efdce36ec8b);
		test(64'ha597eb1117cd8f5a, 64'h1cb2ccae72e282c4, 64'h0000000006f8079a, 64'h14b20c2832a08240, 64'h5a79be1171dcf8a5);
		test(64'hdc42c1092b7d76c1, 64'hc237b2f270761c6c, 64'h00000000c2802f58, 64'h021332d070321004, 64'hd7b21c6724cd901c);
		test(64'h6a0bba3d9c346b54, 64'h3e265f50ca785682, 64'h000000002a5a69a4, 64'h1c00541088681200, 64'h9a0eeac763c19e51);
		test(64'h490020c1727746af, 64'h30a735bd4253e3e2, 64'h000000000110feab, 64'h10a1059c400342e2, 64'hd8dd19af16008034);
		test(64'hae251c6b2919fca5, 64'h5ec624fa0a98461c, 64'h000000000392dcf1, 64'h440600fa08104014, 64'hb6c152ea5acf9192);
		test(64'h35a977dcb37f7190, 64'h9384339fed11eb73, 64'h00000002dfe53b24, 64'h8104218fe5102840, 64'he890dcefeeb3ca59);
		test(64'h569f761f43157465, 64'hf7ae0bc4d9d8e7cd, 64'h000000175d14938b, 64'h76800a0448d08309, 64'hf69af29ba238a98b);
		test(64'h4d074888302f0542, 64'h617ff45c5cb64bc8, 64'h000000050e82458a, 64'h0018105c00244040, 64'h074d88482f304205);
		test(64'hb0a196fcaa5ad55f, 64'h7c1bc191317ad735, 64'h00000000c19a5fd7, 64'h2812409021524535, 64'haefa555a96cf0725);
		test(64'h6cc39ae788fd4fdb, 64'hb5fff7a7964c2384, 64'h0000000ac395f8ee, 64'h1588f68496482284, 64'hc63ca97e88dff4bd);
		test(64'h6d548f557b9edac3, 64'h458a876882eb37b6, 64'h0000000071f19951, 64'h4582846880ca2606, 64'ha7c3edb6f2557915);
		test(64'ha57a47b01767cc59, 64'h57fbf3b43c333581, 64'h00000002be4f96c9, 64'h002b61b40c011401, 64'h5ab58b702b9bcca6);
		test(64'hf46a12b6196213aa, 64'he722777b95bb7d0d, 64'h0000007994d2a44c, 64'h6300145810116904, 64'h598f971219625532);
		test(64'h9710581ab280e8b7, 64'hcd875dc4738524a6, 64'h000000004c381d2f, 64'h4882004450042426, 64'h8e022bded60425a4);
		test(64'h7e54d16c3061c76f, 64'hae2c34f4b6df3f21, 64'h0000000794d6211f, 64'ha00c003006871b21, 64'h3092cb9fbda8e29c);
		test(64'ha635d859dda7691f, 64'h21514be1eaff800d, 64'h00000000278baa77, 64'h01504921a891800d, 64'ha3956a4eb5eef269);
		test(64'h509be1c4de51dc4d, 64'h550fccdd6179ccb5, 64'h000000065e652be3, 64'h410bc09061380831, 64'hcee8de2a2d8c0a76);
		test(64'h3daa308ed886b26c, 64'h43def9e47ac6a408, 64'h00000000329936bd, 64'h42c209444844a000, 64'haa3d8e3086d86cb2);
		test(64'hf9781c67819b2b40, 64'hf0199ff9d716cd16, 64'h0000000fce330d28, 64'h7010033185064000, 64'h34d96f2de80142e6);
		test(64'h12c31903f2b1650c, 64'h32364ac2fc20c4c6, 64'h0000000003147cb2, 64'h10260082940000c0, 64'h84c364c08f4e5930);
		test(64'h68401b8e80ef74cf, 64'h3bef3950bb6679e6, 64'h0000002881c83f9b, 64'h0b400940b9621866, 64'h02fb1df32901e4b2);
		test(64'h95bcbd0415980c95, 64'h0d88f38d09bab9cc, 64'h000000003ed26c29, 64'h0108618000182144, 64'hcb5940db895159c0);
		test(64'h53e0f46355403fbf, 64'hc21bcfd3a412b000, 64'h0000000001868b23, 64'h401001d38412b000, 64'h53e0f46355403fbf);
		test(64'h4ad8dbca7b369560, 64'hfe093616b05da04a, 64'h0000000009652d54, 64'hd809141090150000, 64'h721a3a7ec9de9065);
		test(64'h36c00b65ad48498a, 64'hf8a19dd2ca03fb99, 64'h00000000d0a9425a, 64'h6821144008013088, 64'h9a07c0394586845e);
		test(64'h2cbad32fe4463a2e, 64'h55c24b7396f1fdda, 64'h000000056d748383, 64'h15c241020611a158, 64'h8f7cea838bca19b1);
		test(64'hdf2885eea35a28a1, 64'h3847a023c4e294b0, 64'h0000000000c2d146, 64'h2806800140208010, 64'h28a1a35a85eedf28);
		test(64'h73c68dbe126a7d99, 64'hf9ecdba96526ef22, 64'h0000000ee65e0af4, 64'hf0208a882524c602, 64'h489ad766dc3927eb);
		test(64'heb9b8385f74b2a7c, 64'h4cf07d570d70a328, 64'h000000003482571b, 64'h48e049420910a300, 64'h4bf77c2a9beb8583);
		test(64'h105dff8ffbfb886e, 64'h1f118f36221fa4fe, 64'h000000010fe7ee37, 64'h1f108f32220200dc, 64'hb922efeff2ff7504);
		test(64'h656cdfb9f5436437, 64'h52c1a33fa4880f3f, 64'h00000000457cf137, 64'h52408206a0080037, 64'hec26c2af9dfb36a6);
		test(64'h5068eb4b99e730e1, 64'h7b14b94e5c84e6c0, 64'h000000002837ad93, 64'h311489424004c040, 64'h5068eb4b99e730e1);
		test(64'hfd93f383c3c65f0d, 64'h1b3db0839fd1b0f3, 64'h0000000353fc7841, 64'h1b01b00092d18031, 64'haf0b3c36fc1cfb9c);
		test(64'h9d892dc7c4384f52, 64'hd4952e791ad1ab4c, 64'h00000000b9e8823c, 64'hc010064010d12208, 64'h98d97cd2834c25f4);
		test(64'h03ca6af7dfd35b1a, 64'h3e56e79d59817b2c, 64'h0000000065adff7a, 64'h3e16e50c49014308, 64'h3dfda1b5ac307fa6);
		test(64'hef085e2649bd32da, 64'hf97a964cb047be3f, 64'h0000001d89c8565a, 64'h3048144c9003161a, 64'h5b4cbd92647a10f7);
		test(64'h666df85a72095e83, 64'h2e3aa5a276968cfe, 64'h00000002eb0f41c1, 64'h2230800212168406, 64'hc2b5608da52f7999);
		test(64'h97377a28fa895e67, 64'h7be4c47d48d1351b, 64'h0000000059a53963, 64'h3b44004908d0140b, 64'h41e5ce9e6ea719f5);
		test(64'h95d6fae0c3ccb1b1, 64'ha4a739feae756492, 64'h00000005b7708c96, 64'h00a019988c146002, 64'hfab06579e4e43c33);
		test(64'hf8cf182db754eadb, 64'h6cc8732d8fc795ce, 64'h00000007727dd91d, 64'h4c483224838514c6, 64'hf32f782415dee7ab);
		test(64'h50c93659854ea965, 64'h731563782a2ccd77, 64'h0000000142d61d75, 64'h6004423808240945, 64'h95a6a1726c9a0a93);
		test(64'hfb27033b9abf292d, 64'hfa6fbe47df1bbc3f, 64'h00000fd704ed7aad, 64'h306b8c42de09102d, 64'hb494fd59dcc0e4df);
		test(64'h1be3c8b528c36487, 64'h6cdcbac059c7238e, 64'h000000002c4a2dcb, 64'h088480c01841000e, 64'hcbe45e23c328d219);
		test(64'h8b452100505f8e49, 64'hed808cf6b0ff8315, 64'h00000001280057f1, 64'h240000b6a0390101, 64'h210074a8d4680afa);
		test(64'h315f4264a0ba1953, 64'h3b1ff971b71559a1, 64'h0000000cfd0cc239, 64'h1108295006044821, 64'h507526a332af8198);
		test(64'h9da1d83e4cbd3b52, 64'h1cfe2d8b1348d5a4, 64'h000000007a08c128, 64'h10ca2c8112484420, 64'hc4dbb325d91a8de3);
		test(64'h7a064aa297f1ad0f, 64'hcaec8a45c03eed95, 64'h0000000070b162f3, 64'h826c8a00c0164095, 64'h58155b90e5f0b62f);
		test(64'haf5e494833ab550e, 64'h25fde6d223f08024, 64'h000000001d7213d1, 64'h20e9624202108020, 64'h33ba55e0fae59484);
		test(64'h43c73acebbdbe824, 64'h050a8acb00bad6f4, 64'h0000000002bf5f05, 64'h010a828b00a80220, 64'h8e42bbbda3ec347c);
		test(64'hcee888a8de629e59, 64'h0ec6e1279ef8ed25, 64'h00000003e447d931, 64'h0286c02414782501, 64'hde19d66adc4d4445);
		test(64'h7efd32689924f5bf, 64'h5b1c7e36f8b43394, 64'h00000003dd989aef, 64'h08182410f0941394, 64'h2386e7df5ffb9942);
		test(64'hfdb7681443dd3ef3, 64'h07cafc398b57584e, 64'h0000000165a43eb9, 64'h0100f43103555806, 64'hde7f142977c1cfbc);
		test(64'hf56edbf58c62257e, 64'hbb163c15c6347eb4, 64'h00000001cb6f5127, 64'ha110180102042eb0, 64'h52e7c826bd5f5fe6);
		test(64'h27d8733899e33b49, 64'h1465f02ae9890f7f, 64'h0000000061f4edc9, 64'h1024702060890649, 64'h92dcc7991cce1be4);
		test(64'h73b793adbab422a1, 64'hc1a431894dd5c2a4, 64'h0000000003efa58e, 64'h4084210008448004, 64'hab4b221a377b39da);
		test(64'h231d16d712284021, 64'h7632074b4fda38e1, 64'h000000004ad62103, 64'h0410010804001001, 64'h21148012132e29eb);
		test(64'h866c09c2417794d0, 64'hd5843c7bf5784ff9, 64'h000000249448f134, 64'h01002013b5104340, 64'he068bb82c1069c49);
		test(64'hfa0dfead97326126, 64'hbcf5659254688c64, 64'h000000003c1f4683, 64'h2c94209000408060, 64'h79231662afd0efda);
		test(64'h52e5579ef397c47c, 64'hb01902e33ae674f4, 64'h0000000009cb672f, 64'ha00902213a0414e0, 64'h4cc73f7975e9255e);
		test(64'h4f8cf85481aa051d, 64'h184561a66e25b657, 64'h000000001588104d, 64'h0000608440012055, 64'h1f2af231a0b88155);
		test(64'h2b6d75870ca888fb, 64'hdaa25c2337d8872a, 64'h000000000d6b24c7, 64'h0a0214002108870a, 64'ha203fe22978e2dd5);
		test(64'h7d5f584aee3bbca4, 64'hc477acbe472662dd, 64'h00000003bc85eaa2, 64'h407380b643242088, 64'h584afaeb85c773dd);
		test(64'h78a7d8444cdb3958, 64'h9c51243327f3d92a, 64'h000000003101373a, 64'h8440241224e14900, 64'h7e1352c6add21172);
		test(64'h653f6292ae5f3418, 64'h521019ace2ad8c70, 64'h00000000024459c9, 64'h401009a860800c00, 64'h3418ae5f6292653f);
		test(64'hcc628df93755cb68, 64'hbc6d420cdcd8bafe, 64'h00000004f04569b4, 64'h1065400894c098d0, 64'h29e355dc6f728933);
		test(64'h144d48040c06740b, 64'h1818c413ff441a23, 64'h0000000002500c63, 64'h0000001274000203, 64'h0306e20d822b2102);
		test(64'h1d829b7c7f567ad7, 64'hd30ff4669aa883e2, 64'h00000000294b9c2d, 64'h530ea44298888162, 64'hdf59da7d47286ed3);
		test(64'h6f23faff390b6a65, 64'hdb97343b630d45f1, 64'h0000000171efad8d, 64'hc382002a61040521, 64'h959a3607f5ff9f13);
		test(64'hccbe84a27850033a, 64'h206ccfb173bf2dbc, 64'h00000003c99c202e, 64'h0020cc10400121a8, 64'ha33005872a48ebcc);
		test(64'h10e3e24c62eabce7, 64'h19e914f477a0b05e, 64'h000000004e89cbf3, 64'h182114505700b00e, 64'h318bcb04db3eab89);
		test(64'hd169b7e42c1426be, 64'hd65ed326a7746173, 64'h00000007297cc34e, 64'h804c010402304172, 64'h46d74382de72b869);
		test(64'hebad05ded1eeb571, 64'haf3970c0e9f8145b, 64'h00000000eec79ef9, 64'ha41950c049501441, 64'hb70a5b7de8da77b8);
		test(64'hde6b066f31c392b3, 64'he4f477b25fbed956, 64'h000000d60ca8c345, 64'h60f030b007124906, 64'h90f9b7e986ce4cc3);
		test(64'h1aac27076d553164, 64'h390172e614e34206, 64'h0000000000c51a92, 64'h2801222400a20200, 64'ha43ad8d079554c19);
		test(64'h01461baf025ec502, 64'hfb91ba85e35b7808, 64'h00000000041f8bd0, 64'h80809a8181100800, 64'h4601af1b5e0202c5);
		test(64'hc49e2666c8b2ccf8, 64'hb54eba915ecd9761, 64'h000000049d2290a6, 64'ha50412804c489700, 64'hc471ccf4c86d1999);
		test(64'h320c539995e7f40f, 64'h86c1dc8691fed827, 64'h000000002193f3e7, 64'h80815c0291e80027, 64'ha9e72ff04c30ca99);
		test(64'he563dc7ba0c1cc57, 64'h7db7cdc02a67ba0f, 64'h0000000cd3f32327, 64'h5c80c0002a061207, 64'hc6a7de3b8305ea33);
		test(64'h2b3c5e25e9ea16bb, 64'h8404260882c70c56, 64'h000000000002d695, 64'h8004000080c20c46, 64'hb558e83c94ee6bab);
		test(64'h78bd3b2a6c1757ce, 64'h52ec698342214ae1, 64'h00000000035dd4dc, 64'h00246102422140e0, 64'h9c2babcdb47e3715);
		test(64'hadea7293c5c39034, 64'h1600bb6ad4829a14, 64'h00000000009a1df3, 64'h1600034200009200, 64'h2739daae09435c3c);
		test(64'h751ddfa6468f9a20, 64'h45c6701940880d14, 64'h00000000001ca8f0, 64'h05c4300800080000, 64'hfd6a57d1a90264f8);
		test(64'h2fa271e9e1b4d80e, 64'h87d5fbc4203c723e, 64'h00000000f073bb47, 64'h8701b2440030001c, 64'hb0271e4b6b4d8af8);
		test(64'h72a47772a393455a, 64'h933f221a200e7550, 64'h0000000001a4eccf, 64'h9213020020045440, 64'h777272a4455aa393);
		test(64'h4a3d2c25a20d3dba, 64'h38cf7036df330941, 64'h000000001355421c, 64'h100810245d230840, 64'h853e1c1a510e3e75);
		test(64'ha66a064921411f13, 64'h2f25e569b37c39ed, 64'h0000001682b4c1c1, 64'h09010120021c3045, 64'h282132f259956890);
		test(64'h17efb2f20d951ade, 64'hc13ecf80a145476b, 64'h000000000de29656, 64'h012c45000141066a, 64'h9a0bb7857f8ef4d4);
		test(64'h94c1f569b7f17725, 64'h9f19765f4f31fc8b, 64'h000000343ea4fdd1, 64'h8911565c0b21c809, 64'h389269faf8de4aee);
		test(64'hc5bd3e05b925ddb2, 64'h86dff31e3584ba89, 64'h000000035d38b5b4, 64'h0659210e15049808, 64'h7eca0a3d1a7671ee);
		test(64'he3c6b2e59ce831bc, 64'h5f05e2ae76540edf, 64'h0000000475e8d05c, 64'h4c0582a40240065c, 64'ha74d63c73d8c1739);
		test(64'hfaeef0fddc64f102, 64'h7777e867d0003860, 64'h000000001d6dddf8, 64'h7062684100000040, 64'hdc64f102faeef0fd);
		test(64'h43e9d50758822010, 64'h216dc91972192050, 64'h00000000007ba685, 64'h2001010000080000, 64'hd50743e920105882);
		test(64'h6c57bfeaee9f0610, 64'hf5674f7e0479bc1c, 64'h00000006aefd670c, 64'ha547097800180800, 64'haefb75c60160f9ee);
		test(64'h216c3dd54155c864, 64'hd6333787f241faf4, 64'h0000000047751e4d, 64'h4420050570010a20, 64'h8c461455d35d12c6);
		test(64'h2d1aeb56da874401, 64'hd05caca0ebf16ac9, 64'h000000000dc6d181, 64'hc0542000e2200001, 64'h251ea9d74be50288);
		test(64'h0439d6f74f9d1a5c, 64'hdc6f3b648bdf3768, 64'h00000002cabbdd55, 64'hcc493a24821a1340, 64'h9d4f5c1a3904f7d6);
		test(64'h61e30a9bf5e45306, 64'h292f7638053b9a20, 64'h000000000b30be0a, 64'h082e202800300a00, 64'hf5e4530661e30a9b);
		test(64'h8a83375482bb6514, 64'h052aa7c64479d6de, 64'h000000000bd87a8a, 64'h040022c444309048, 64'h15dcc2a21459ee82);
		test(64'hc65e132949b952f3, 64'h9ce7f22ba60cfc96, 64'h00000004ac3d094d, 64'h0884d2212200bc06, 64'hc46893b585cf616e);
		test(64'he5a8183dec3300ef, 64'h12830c9d816abd2e, 64'h00000000024f940f, 64'h1200048500001c2e, 64'hcc3bfb002a5b7c24);
		test(64'h4865f30c70cae3d4, 64'h1c36783d00cf0313, 64'h0000000002ae375c, 64'h00305038004e0210, 64'hfc03216a7cb2e035);
		test(64'ha5bee94cdac639d5, 64'hc186377ef40b60e6, 64'h00000000be33693a, 64'hc0842618700340a2, 64'ha7936c575abe6b31);
		test(64'h733ff46378698fa7, 64'h7419d6443ffe5578, 64'h000000077f5c3434, 64'h30198044131e4438, 64'ha78f697863f43f73);
		test(64'ha87df66f6d1ff7d2, 64'he16b6e7ff3b87cbd, 64'h000002bbbdec9f68, 64'h814b4c68f3b07c24, 64'h1ebff2e9f99feb45);
		test(64'h3fec0287ebdf8304, 64'hb2c44113198c7d02, 64'h0000000000fc6f82, 64'hb0c4411000880400, 64'hcfb3082dbe7f2c01);
		test(64'he65e486619f06578, 64'h739164a51211dbb2, 64'h000000001a51a916, 64'h6191400110014b80, 64'h95d246f01299b95b);
		test(64'hc56e03004e3f5485, 64'h28a0411f7d3eab6c, 64'h000000000a09be01, 64'h2020410379142024, 64'hf3e45845e65c0030);
		test(64'h73091be2c3778d3a, 64'h02c3fc61f3f56ca0, 64'h0000000088db37cd, 64'h02806c41e0d06880, 64'hc3778d3a73091be2);
		test(64'hc6839c203c2fae79, 64'h9d4890741cb94f65, 64'h000000002469d6ed, 64'h9c00103418990741, 64'hc3f1d56b9c34c601);
		test(64'hb1d179ba7a4944bb, 64'h6ae69269859f98f2, 64'h00000000984c0917, 64'h0ac41020810488d2, 64'h11eeda16d6eae474);
		test(64'h52e5714674eadb43, 64'hb47d171fe5b7be35, 64'h0000002ce4cecad1, 64'h2031150744a6a805, 64'h7e388b5d2b981aad);
		test(64'hba4f56d5b847fc09, 64'hc409308c5e2b51b1, 64'h00000000026d61e1, 64'h0008008c5e200081, 64'hfc06748ba9ea758f);
		test(64'hf7a3c6d530d14b52, 64'haa7a9d1e7d007d44, 64'h00000000d4ca9896, 64'h0a02880a15002840, 64'h7f3a6c5d031db425);
		test(64'h381cfc805731acbe, 64'h79d6b34ceead2067, 64'h000000038dc09a6e, 64'h01468300ca842066, 64'hea8c357d1c383f01);
		test(64'h0f68a0ad7ffa83e7, 64'hf1d2e2fe55996f20, 64'h0000000052ab7f07, 64'ha1d2e2ea00196320, 64'h7ffa83e70f68a0ad);
		test(64'hc8edf706c97195fe, 64'h1e0860073893c955, 64'h00000000009f159e, 64'h160800030811c954, 64'hbf904ceda6df6c2b);
		test(64'h3e1a406f5c341b87, 64'h7f879d4ae81a7270, 64'h00000000f881d618, 64'h57009400601a0070, 64'h1b875c34406f3e1a);
		test(64'hb6a4f7f88030da94, 64'h88699c985a169e21, 64'h00000000049bc274, 64'h0001801818120a00, 64'h4030e5687958fbf4);
		test(64'h7f671b770a7b1b5d, 64'h4ea9da492d949a2b, 64'h000000007a9ea275, 64'h0220d84805141229, 64'hed05ab8d6eefee8d);
		test(64'h0903ad5cfa1259df, 64'hb8a47aed5913eaac, 64'h000000004296ecab, 64'h18a420441110e2ac, 64'h21affd953090c5da);
		test(64'h734f567176fce679, 64'h6c0d1590f40da1f5, 64'h0000000019f2fd9d, 64'h4c051580700501e1, 64'h9d6b9bcf9a2b3bf8);
		test(64'h252cb061ad5f67f6, 64'h3bc56e841c50e4b9, 64'h0000000022481efc, 64'h2a846e041050e498, 64'hf99baf5e92701c1a);
		test(64'h1a91ff588aa64b30, 64'h1290ad5fcc0bcba6, 64'h000000007ff8a4f4, 64'h0010244640098300, 64'ha29ae10ca446ff25);
		test(64'h43db325ce377f5b1, 64'h3b077c9ad5ce561a, 64'h000000006d8d95f4, 64'h0b006c8ad5461402, 64'h53c87e1ce4f5ddbc);
		test(64'hc9e3bc09415f0c36, 64'h1d0b9a3a1ac47fae, 64'h00000000af88318b, 64'h1400121a1800618c, 64'hf5419c30cb63603e);
		test(64'hef30e0e7e9b9dcd1, 64'h791ca2e405d7bb28, 64'h000000006e6f69b0, 64'h680c22840554a808, 64'hb9e9d1dc30efe7e0);
		test(64'ha8ae3cb5f3ebde5e, 64'h887cc1ada5f45e62, 64'h00000000d637bcfd, 64'h8864c189a4f01660, 64'hfcbe7b5ba2abc3e5);
		test(64'hdf9bf731d4d86e5e, 64'hcc5c2f729ea58902, 64'h000000003daeda85, 64'h440c0c121c218900, 64'h7f6efdc471729b5b);
		test(64'h799fdfeae6fac290, 64'h0f01ed98f3ff9315, 64'h00000004f7bd7d54, 64'h05018c98d1850200, 64'hfe5d6bf61c069d5f);
		test(64'h1ed6093cdd780973, 64'h3d23866b70acc5a1, 64'h000000001c832b0b, 64'h1c2186001008c421, 64'heeb406b32de9063c);
		test(64'h26291e3fbd1cd46a, 64'h6d7b0bf2715ab742, 64'h0000000295c776b3, 64'h6c7900e061103240, 64'h89864bcfe743719a);
		test(64'h92b864a9b0a592ac, 64'h8f21f9f39de7f289, 64'h00000025314e2d9e, 64'h842160508c42a280, 64'h746156985a705c61);
		test(64'hdbc84fb88329bf2c, 64'h915f3e294101a752, 64'h000000000f41f3f8, 64'h01450c2941010540, 64'h1fe27e32ef832c86);
		test(64'h323dec250638309c, 64'hf251b62c0bd1e7fd, 64'h00000003bd54444e, 64'h5000300c08018138, 64'hc6034390a1cde313);
		test(64'hfb6c29b8ada41b72, 64'h6a4fe75ba91fcfc4, 64'h0000003f84b3c85a, 64'h68056311000d8e40, 64'hbfc6928bda4ab127);
		test(64'h21309bd1a2f0815b, 64'h478f61ac008c5699, 64'h000000000080c407, 64'h058c010000041289, 64'he2673012a742f051);
		test(64'h821076e961a3c874, 64'h0d058550875412e4, 64'h0000000000014207, 64'h0400854004041240, 64'h163a8c472801679e);
		test(64'h29f62894768083c1, 64'h332cb3624b395286, 64'h000000001350280c, 64'h2308002000390002, 64'h689f28169d02c243);
		test(64'h53e8aca7e8ed41a3, 64'h14c2c1a8139893e0, 64'h0000000000b4c28d, 64'h1482812000181060, 64'he8ed41a353e8aca7);
		test(64'h14d7439202695ac7, 64'h6eed671f2407d9b2, 64'h00000000b39c82e9, 64'h2004250504055032, 64'h5a3d08961c68417d);
		test(64'hfebb5f87158dfa81, 64'hc0f8a55c05e06134, 64'h0000000003b98f30, 64'h4088855c01400004, 64'haf1851d8f578efbb);
		test(64'hd2ac100110396cf6, 64'h84c909dbf682e3af, 64'h0000000150088336, 64'h8008000b260283a6, 64'h9c086f36354b8008);
		test(64'h8372e8a066f2eda8, 64'h8cb7a7d403d76273, 64'h000000023588bac8, 64'h00a3271003954220, 64'h7b5166f471501ce4);
		test(64'h037ed96dd2a83077, 64'h521e8fe19ea19dd7, 64'h00000001fcbe721f, 64'h421a054100a001c7, 64'h9bb6c07e0cee4b15);
		test(64'h707ef5cf50194b2c, 64'h8c7d52ef84fa32ba, 64'h00000000fb6f062a, 64'h8c280029042a0230, 64'h831e46503ff5dbd0);
		test(64'he004a5647396285f, 64'h82c04ca17c6ef3cf, 64'h0000000082b8321f, 64'h02c004a02c04814f, 64'h200726a569cefa14);
		test(64'h1d973d4c80833de8, 64'h5bc66de6ddd64193, 64'h00000006dbd50458, 64'h510004028d964080, 64'hcb238b9ecb71101c);
		test(64'h113718af7e6fe9d0, 64'h96de3e2ac2554203, 64'h00000000085b3bb8, 64'h961a3e2202510000, 64'h88ce815fe76f79b0);
		test(64'hf0e0052eba4f0847, 64'h422272215adf6797, 64'h00000000504ebc07, 64'h022220201a820207, 64'ha0740f0710e25df2);
		test(64'h27ee134bfa71dc98, 64'h21f7f61ff8231921, 64'h00000001f6157fb8, 64'h21f2700ee0201800, 64'hf5b2ec641bdd2387);
		test(64'h1c99396bc2973753, 64'h68b585d00dcfadfd, 64'h00000001a94275a9, 64'h28a0048009c32ca5, 64'h3ab3b61c796366c2);
		test(64'hef7dcc60f04cede6, 64'h35c74f9a2451cdbd, 64'h00000002dbc0a7f2, 64'h05c0049024418d8c, 64'h9dedc80f09ccebfd);
		test(64'h1b8018bd7f11a166, 64'h28c57367c2e31ba4, 64'h000000003046b08b, 64'h28c54103400218a0, 64'hf7111a66b10881db);
		test(64'h37ff7584bff2b493, 64'h238144da36c6153a, 64'h0000000007f87ee5, 64'h238144121482010a, 64'h6ce1f8ef21d5ffcd);
		test(64'h6701d515dea99790, 64'h0d22f31b2cfd20bf, 64'h00000000cd65d550, 64'h0d02e2120c2d2010, 64'h09e9957ba8ab80e6);
		test(64'h78b4165fab87153e, 64'hc259338c3e9a9494, 64'h000000000919d65b, 64'h405801880a109490, 64'h61f5874b51e3ba78);

		@(posedge clk);
		$display("Final cycle count: %1d", cycles);
		$display("OK");
		$finish;
	end
endmodule
