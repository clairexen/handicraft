
`include "common.svh"

module top();
  type_fruit_e fruit;
  mymodule uut(
      .fruit(fruit)
  );
endmodule

