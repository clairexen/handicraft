
module regcell(
	\input , enable, Q
);

input [2:0] \input ;
input enable;
output [2:0] Q;

/* leave the module empty - xst will recognice it as blackbox module */

endmodule

