
`include "common.svh"

module mymodule(output type_fruit_e fruit);
    assign fruit = APPLE;
endmodule
