`timescale 1ns / 1ps
module PROM(
    input [10:0] adr,
    output reg [31:0] data,
    input clk);
reg [31:0] mem [2047: 0];
initial $readmemh("prom.mem", mem);
always @(posedge clk) data <= mem[adr];
endmodule

