module top(input A, output Y);
  assign Y = !A;
endmodule
