module testbox_A(input A, B, output Y);
assign Y = A;
endmodule
