
typedef enum logic[1:0] {
    APPLE               = 2'b00,
    BANANA              = 2'b01,
    ORANGE              = 2'b10,
    PEAR                = 2'b11
} type_fruit_e;

