module testbox_B(input A, B, output Y);
assign Y = B;
endmodule
