module dummy (input in, output out);
  assign out = in;
endmodule
